module heichips25_SDR (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.I_range.data_plus_4[6] ;
 wire \DP_1.I_range.out_data[2] ;
 wire \DP_1.I_range.out_data[3] ;
 wire \DP_1.I_range.out_data[4] ;
 wire \DP_1.I_range.out_data[5] ;
 wire \DP_1.I_range.out_data[6] ;
 wire \DP_1.Q_range.data_plus_4[6] ;
 wire \DP_1.Q_range.out_data[2] ;
 wire \DP_1.Q_range.out_data[3] ;
 wire \DP_1.Q_range.out_data[4] ;
 wire \DP_1.Q_range.out_data[5] ;
 wire \DP_1.Q_range.out_data[6] ;
 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[2] ;
 wire \DP_1.matrix[36] ;
 wire \DP_1.matrix[37] ;
 wire \DP_1.matrix[38] ;
 wire \DP_1.matrix[39] ;
 wire \DP_1.matrix[3] ;
 wire \DP_1.matrix[40] ;
 wire \DP_1.matrix[41] ;
 wire \DP_1.matrix[42] ;
 wire \DP_1.matrix[43] ;
 wire \DP_1.matrix[44] ;
 wire \DP_1.matrix[4] ;
 wire \DP_1.matrix[5] ;
 wire \DP_1.matrix[6] ;
 wire \DP_1.matrix[72] ;
 wire \DP_1.matrix[73] ;
 wire \DP_1.matrix[74] ;
 wire \DP_1.matrix[75] ;
 wire \DP_1.matrix[76] ;
 wire \DP_1.matrix[77] ;
 wire \DP_1.matrix[78] ;
 wire \DP_1.matrix[79] ;
 wire \DP_1.matrix[7] ;
 wire \DP_1.matrix[80] ;
 wire \DP_1.matrix[8] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[2] ;
 wire \DP_2.matrix[36] ;
 wire \DP_2.matrix[37] ;
 wire \DP_2.matrix[38] ;
 wire \DP_2.matrix[39] ;
 wire \DP_2.matrix[3] ;
 wire \DP_2.matrix[40] ;
 wire \DP_2.matrix[41] ;
 wire \DP_2.matrix[42] ;
 wire \DP_2.matrix[43] ;
 wire \DP_2.matrix[44] ;
 wire \DP_2.matrix[4] ;
 wire \DP_2.matrix[5] ;
 wire \DP_2.matrix[6] ;
 wire \DP_2.matrix[72] ;
 wire \DP_2.matrix[73] ;
 wire \DP_2.matrix[74] ;
 wire \DP_2.matrix[75] ;
 wire \DP_2.matrix[76] ;
 wire \DP_2.matrix[77] ;
 wire \DP_2.matrix[78] ;
 wire \DP_2.matrix[79] ;
 wire \DP_2.matrix[7] ;
 wire \DP_2.matrix[80] ;
 wire \DP_2.matrix[8] ;
 wire \DP_3.I_range.data_plus_4[6] ;
 wire \DP_3.I_range.out_data[2] ;
 wire \DP_3.I_range.out_data[3] ;
 wire \DP_3.I_range.out_data[4] ;
 wire \DP_3.I_range.out_data[5] ;
 wire \DP_3.I_range.out_data[6] ;
 wire \DP_3.Q_range.data_plus_4[6] ;
 wire \DP_3.Q_range.out_data[2] ;
 wire \DP_3.Q_range.out_data[3] ;
 wire \DP_3.Q_range.out_data[4] ;
 wire \DP_3.Q_range.out_data[5] ;
 wire \DP_3.Q_range.out_data[6] ;
 wire \DP_3.matrix[0] ;
 wire \DP_3.matrix[1] ;
 wire \DP_3.matrix[2] ;
 wire \DP_3.matrix[36] ;
 wire \DP_3.matrix[37] ;
 wire \DP_3.matrix[38] ;
 wire \DP_3.matrix[39] ;
 wire \DP_3.matrix[3] ;
 wire \DP_3.matrix[40] ;
 wire \DP_3.matrix[41] ;
 wire \DP_3.matrix[42] ;
 wire \DP_3.matrix[43] ;
 wire \DP_3.matrix[44] ;
 wire \DP_3.matrix[4] ;
 wire \DP_3.matrix[5] ;
 wire \DP_3.matrix[6] ;
 wire \DP_3.matrix[72] ;
 wire \DP_3.matrix[73] ;
 wire \DP_3.matrix[74] ;
 wire \DP_3.matrix[75] ;
 wire \DP_3.matrix[76] ;
 wire \DP_3.matrix[77] ;
 wire \DP_3.matrix[78] ;
 wire \DP_3.matrix[79] ;
 wire \DP_3.matrix[7] ;
 wire \DP_3.matrix[80] ;
 wire \DP_3.matrix[8] ;
 wire \DP_4.matrix[0] ;
 wire \DP_4.matrix[1] ;
 wire \DP_4.matrix[2] ;
 wire \DP_4.matrix[36] ;
 wire \DP_4.matrix[37] ;
 wire \DP_4.matrix[38] ;
 wire \DP_4.matrix[39] ;
 wire \DP_4.matrix[3] ;
 wire \DP_4.matrix[40] ;
 wire \DP_4.matrix[41] ;
 wire \DP_4.matrix[42] ;
 wire \DP_4.matrix[43] ;
 wire \DP_4.matrix[44] ;
 wire \DP_4.matrix[4] ;
 wire \DP_4.matrix[5] ;
 wire \DP_4.matrix[6] ;
 wire \DP_4.matrix[72] ;
 wire \DP_4.matrix[73] ;
 wire \DP_4.matrix[74] ;
 wire \DP_4.matrix[75] ;
 wire \DP_4.matrix[76] ;
 wire \DP_4.matrix[77] ;
 wire \DP_4.matrix[78] ;
 wire \DP_4.matrix[79] ;
 wire \DP_4.matrix[7] ;
 wire \DP_4.matrix[80] ;
 wire \DP_4.matrix[8] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[10] ;
 wire \mac1.products_ff[11] ;
 wire \mac1.products_ff[12] ;
 wire \mac1.products_ff[136] ;
 wire \mac1.products_ff[137] ;
 wire \mac1.products_ff[138] ;
 wire \mac1.products_ff[139] ;
 wire \mac1.products_ff[13] ;
 wire \mac1.products_ff[140] ;
 wire \mac1.products_ff[141] ;
 wire \mac1.products_ff[142] ;
 wire \mac1.products_ff[143] ;
 wire \mac1.products_ff[144] ;
 wire \mac1.products_ff[145] ;
 wire \mac1.products_ff[146] ;
 wire \mac1.products_ff[147] ;
 wire \mac1.products_ff[148] ;
 wire \mac1.products_ff[149] ;
 wire \mac1.products_ff[14] ;
 wire \mac1.products_ff[150] ;
 wire \mac1.products_ff[151] ;
 wire \mac1.products_ff[15] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[2] ;
 wire \mac1.products_ff[3] ;
 wire \mac1.products_ff[4] ;
 wire \mac1.products_ff[5] ;
 wire \mac1.products_ff[68] ;
 wire \mac1.products_ff[69] ;
 wire \mac1.products_ff[6] ;
 wire \mac1.products_ff[70] ;
 wire \mac1.products_ff[71] ;
 wire \mac1.products_ff[72] ;
 wire \mac1.products_ff[73] ;
 wire \mac1.products_ff[74] ;
 wire \mac1.products_ff[75] ;
 wire \mac1.products_ff[76] ;
 wire \mac1.products_ff[77] ;
 wire \mac1.products_ff[78] ;
 wire \mac1.products_ff[79] ;
 wire \mac1.products_ff[7] ;
 wire \mac1.products_ff[80] ;
 wire \mac1.products_ff[81] ;
 wire \mac1.products_ff[82] ;
 wire \mac1.products_ff[83] ;
 wire \mac1.products_ff[8] ;
 wire \mac1.products_ff[9] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[10] ;
 wire \mac1.sum_lvl1_ff[11] ;
 wire \mac1.sum_lvl1_ff[12] ;
 wire \mac1.sum_lvl1_ff[13] ;
 wire \mac1.sum_lvl1_ff[14] ;
 wire \mac1.sum_lvl1_ff[15] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[2] ;
 wire \mac1.sum_lvl1_ff[36] ;
 wire \mac1.sum_lvl1_ff[37] ;
 wire \mac1.sum_lvl1_ff[38] ;
 wire \mac1.sum_lvl1_ff[39] ;
 wire \mac1.sum_lvl1_ff[3] ;
 wire \mac1.sum_lvl1_ff[40] ;
 wire \mac1.sum_lvl1_ff[41] ;
 wire \mac1.sum_lvl1_ff[42] ;
 wire \mac1.sum_lvl1_ff[43] ;
 wire \mac1.sum_lvl1_ff[44] ;
 wire \mac1.sum_lvl1_ff[45] ;
 wire \mac1.sum_lvl1_ff[46] ;
 wire \mac1.sum_lvl1_ff[47] ;
 wire \mac1.sum_lvl1_ff[48] ;
 wire \mac1.sum_lvl1_ff[49] ;
 wire \mac1.sum_lvl1_ff[4] ;
 wire \mac1.sum_lvl1_ff[50] ;
 wire \mac1.sum_lvl1_ff[51] ;
 wire \mac1.sum_lvl1_ff[5] ;
 wire \mac1.sum_lvl1_ff[6] ;
 wire \mac1.sum_lvl1_ff[72] ;
 wire \mac1.sum_lvl1_ff[73] ;
 wire \mac1.sum_lvl1_ff[74] ;
 wire \mac1.sum_lvl1_ff[75] ;
 wire \mac1.sum_lvl1_ff[76] ;
 wire \mac1.sum_lvl1_ff[77] ;
 wire \mac1.sum_lvl1_ff[78] ;
 wire \mac1.sum_lvl1_ff[79] ;
 wire \mac1.sum_lvl1_ff[7] ;
 wire \mac1.sum_lvl1_ff[80] ;
 wire \mac1.sum_lvl1_ff[81] ;
 wire \mac1.sum_lvl1_ff[82] ;
 wire \mac1.sum_lvl1_ff[83] ;
 wire \mac1.sum_lvl1_ff[84] ;
 wire \mac1.sum_lvl1_ff[85] ;
 wire \mac1.sum_lvl1_ff[86] ;
 wire \mac1.sum_lvl1_ff[87] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[10] ;
 wire \mac1.sum_lvl2_ff[11] ;
 wire \mac1.sum_lvl2_ff[12] ;
 wire \mac1.sum_lvl2_ff[13] ;
 wire \mac1.sum_lvl2_ff[14] ;
 wire \mac1.sum_lvl2_ff[15] ;
 wire \mac1.sum_lvl2_ff[19] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[20] ;
 wire \mac1.sum_lvl2_ff[21] ;
 wire \mac1.sum_lvl2_ff[22] ;
 wire \mac1.sum_lvl2_ff[23] ;
 wire \mac1.sum_lvl2_ff[24] ;
 wire \mac1.sum_lvl2_ff[25] ;
 wire \mac1.sum_lvl2_ff[26] ;
 wire \mac1.sum_lvl2_ff[27] ;
 wire \mac1.sum_lvl2_ff[28] ;
 wire \mac1.sum_lvl2_ff[29] ;
 wire \mac1.sum_lvl2_ff[2] ;
 wire \mac1.sum_lvl2_ff[30] ;
 wire \mac1.sum_lvl2_ff[31] ;
 wire \mac1.sum_lvl2_ff[32] ;
 wire \mac1.sum_lvl2_ff[33] ;
 wire \mac1.sum_lvl2_ff[34] ;
 wire \mac1.sum_lvl2_ff[38] ;
 wire \mac1.sum_lvl2_ff[39] ;
 wire \mac1.sum_lvl2_ff[3] ;
 wire \mac1.sum_lvl2_ff[40] ;
 wire \mac1.sum_lvl2_ff[41] ;
 wire \mac1.sum_lvl2_ff[42] ;
 wire \mac1.sum_lvl2_ff[43] ;
 wire \mac1.sum_lvl2_ff[44] ;
 wire \mac1.sum_lvl2_ff[45] ;
 wire \mac1.sum_lvl2_ff[46] ;
 wire \mac1.sum_lvl2_ff[47] ;
 wire \mac1.sum_lvl2_ff[48] ;
 wire \mac1.sum_lvl2_ff[49] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[50] ;
 wire \mac1.sum_lvl2_ff[51] ;
 wire \mac1.sum_lvl2_ff[52] ;
 wire \mac1.sum_lvl2_ff[53] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[6] ;
 wire \mac1.sum_lvl2_ff[7] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[10] ;
 wire \mac1.sum_lvl3_ff[11] ;
 wire \mac1.sum_lvl3_ff[12] ;
 wire \mac1.sum_lvl3_ff[13] ;
 wire \mac1.sum_lvl3_ff[14] ;
 wire \mac1.sum_lvl3_ff[15] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[20] ;
 wire \mac1.sum_lvl3_ff[21] ;
 wire \mac1.sum_lvl3_ff[22] ;
 wire \mac1.sum_lvl3_ff[23] ;
 wire \mac1.sum_lvl3_ff[24] ;
 wire \mac1.sum_lvl3_ff[25] ;
 wire \mac1.sum_lvl3_ff[26] ;
 wire \mac1.sum_lvl3_ff[27] ;
 wire \mac1.sum_lvl3_ff[28] ;
 wire \mac1.sum_lvl3_ff[29] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[30] ;
 wire \mac1.sum_lvl3_ff[31] ;
 wire \mac1.sum_lvl3_ff[32] ;
 wire \mac1.sum_lvl3_ff[33] ;
 wire \mac1.sum_lvl3_ff[34] ;
 wire \mac1.sum_lvl3_ff[35] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.sum_lvl3_ff[4] ;
 wire \mac1.sum_lvl3_ff[5] ;
 wire \mac1.sum_lvl3_ff[6] ;
 wire \mac1.sum_lvl3_ff[7] ;
 wire \mac1.sum_lvl3_ff[8] ;
 wire \mac1.sum_lvl3_ff[9] ;
 wire \mac1.total_sum[0] ;
 wire \mac1.total_sum[10] ;
 wire \mac1.total_sum[11] ;
 wire \mac1.total_sum[12] ;
 wire \mac1.total_sum[13] ;
 wire \mac1.total_sum[14] ;
 wire \mac1.total_sum[15] ;
 wire \mac1.total_sum[1] ;
 wire \mac1.total_sum[2] ;
 wire \mac1.total_sum[3] ;
 wire \mac1.total_sum[4] ;
 wire \mac1.total_sum[5] ;
 wire \mac1.total_sum[6] ;
 wire \mac1.total_sum[7] ;
 wire \mac1.total_sum[8] ;
 wire \mac1.total_sum[9] ;
 wire \mac2.products_ff[0] ;
 wire \mac2.products_ff[10] ;
 wire \mac2.products_ff[11] ;
 wire \mac2.products_ff[12] ;
 wire \mac2.products_ff[136] ;
 wire \mac2.products_ff[137] ;
 wire \mac2.products_ff[138] ;
 wire \mac2.products_ff[139] ;
 wire \mac2.products_ff[13] ;
 wire \mac2.products_ff[140] ;
 wire \mac2.products_ff[141] ;
 wire \mac2.products_ff[142] ;
 wire \mac2.products_ff[143] ;
 wire \mac2.products_ff[144] ;
 wire \mac2.products_ff[145] ;
 wire \mac2.products_ff[146] ;
 wire \mac2.products_ff[147] ;
 wire \mac2.products_ff[148] ;
 wire \mac2.products_ff[149] ;
 wire \mac2.products_ff[14] ;
 wire \mac2.products_ff[150] ;
 wire \mac2.products_ff[151] ;
 wire \mac2.products_ff[15] ;
 wire \mac2.products_ff[1] ;
 wire \mac2.products_ff[2] ;
 wire \mac2.products_ff[3] ;
 wire \mac2.products_ff[4] ;
 wire \mac2.products_ff[5] ;
 wire \mac2.products_ff[68] ;
 wire \mac2.products_ff[69] ;
 wire \mac2.products_ff[6] ;
 wire \mac2.products_ff[70] ;
 wire \mac2.products_ff[71] ;
 wire \mac2.products_ff[72] ;
 wire \mac2.products_ff[73] ;
 wire \mac2.products_ff[74] ;
 wire \mac2.products_ff[75] ;
 wire \mac2.products_ff[76] ;
 wire \mac2.products_ff[77] ;
 wire \mac2.products_ff[78] ;
 wire \mac2.products_ff[79] ;
 wire \mac2.products_ff[7] ;
 wire \mac2.products_ff[80] ;
 wire \mac2.products_ff[81] ;
 wire \mac2.products_ff[82] ;
 wire \mac2.products_ff[83] ;
 wire \mac2.products_ff[8] ;
 wire \mac2.products_ff[9] ;
 wire \mac2.sum_lvl1_ff[0] ;
 wire \mac2.sum_lvl1_ff[10] ;
 wire \mac2.sum_lvl1_ff[11] ;
 wire \mac2.sum_lvl1_ff[12] ;
 wire \mac2.sum_lvl1_ff[13] ;
 wire \mac2.sum_lvl1_ff[14] ;
 wire \mac2.sum_lvl1_ff[15] ;
 wire \mac2.sum_lvl1_ff[1] ;
 wire \mac2.sum_lvl1_ff[2] ;
 wire \mac2.sum_lvl1_ff[36] ;
 wire \mac2.sum_lvl1_ff[37] ;
 wire \mac2.sum_lvl1_ff[38] ;
 wire \mac2.sum_lvl1_ff[39] ;
 wire \mac2.sum_lvl1_ff[3] ;
 wire \mac2.sum_lvl1_ff[40] ;
 wire \mac2.sum_lvl1_ff[41] ;
 wire \mac2.sum_lvl1_ff[42] ;
 wire \mac2.sum_lvl1_ff[43] ;
 wire \mac2.sum_lvl1_ff[44] ;
 wire \mac2.sum_lvl1_ff[45] ;
 wire \mac2.sum_lvl1_ff[46] ;
 wire \mac2.sum_lvl1_ff[47] ;
 wire \mac2.sum_lvl1_ff[48] ;
 wire \mac2.sum_lvl1_ff[49] ;
 wire \mac2.sum_lvl1_ff[4] ;
 wire \mac2.sum_lvl1_ff[50] ;
 wire \mac2.sum_lvl1_ff[51] ;
 wire \mac2.sum_lvl1_ff[5] ;
 wire \mac2.sum_lvl1_ff[6] ;
 wire \mac2.sum_lvl1_ff[72] ;
 wire \mac2.sum_lvl1_ff[73] ;
 wire \mac2.sum_lvl1_ff[74] ;
 wire \mac2.sum_lvl1_ff[75] ;
 wire \mac2.sum_lvl1_ff[76] ;
 wire \mac2.sum_lvl1_ff[77] ;
 wire \mac2.sum_lvl1_ff[78] ;
 wire \mac2.sum_lvl1_ff[79] ;
 wire \mac2.sum_lvl1_ff[7] ;
 wire \mac2.sum_lvl1_ff[80] ;
 wire \mac2.sum_lvl1_ff[81] ;
 wire \mac2.sum_lvl1_ff[82] ;
 wire \mac2.sum_lvl1_ff[83] ;
 wire \mac2.sum_lvl1_ff[84] ;
 wire \mac2.sum_lvl1_ff[85] ;
 wire \mac2.sum_lvl1_ff[86] ;
 wire \mac2.sum_lvl1_ff[87] ;
 wire \mac2.sum_lvl1_ff[8] ;
 wire \mac2.sum_lvl1_ff[9] ;
 wire \mac2.sum_lvl2_ff[0] ;
 wire \mac2.sum_lvl2_ff[10] ;
 wire \mac2.sum_lvl2_ff[11] ;
 wire \mac2.sum_lvl2_ff[12] ;
 wire \mac2.sum_lvl2_ff[13] ;
 wire \mac2.sum_lvl2_ff[14] ;
 wire \mac2.sum_lvl2_ff[15] ;
 wire \mac2.sum_lvl2_ff[19] ;
 wire \mac2.sum_lvl2_ff[1] ;
 wire \mac2.sum_lvl2_ff[20] ;
 wire \mac2.sum_lvl2_ff[21] ;
 wire \mac2.sum_lvl2_ff[22] ;
 wire \mac2.sum_lvl2_ff[23] ;
 wire \mac2.sum_lvl2_ff[24] ;
 wire \mac2.sum_lvl2_ff[25] ;
 wire \mac2.sum_lvl2_ff[26] ;
 wire \mac2.sum_lvl2_ff[27] ;
 wire \mac2.sum_lvl2_ff[28] ;
 wire \mac2.sum_lvl2_ff[29] ;
 wire \mac2.sum_lvl2_ff[2] ;
 wire \mac2.sum_lvl2_ff[30] ;
 wire \mac2.sum_lvl2_ff[31] ;
 wire \mac2.sum_lvl2_ff[32] ;
 wire \mac2.sum_lvl2_ff[33] ;
 wire \mac2.sum_lvl2_ff[34] ;
 wire \mac2.sum_lvl2_ff[38] ;
 wire \mac2.sum_lvl2_ff[39] ;
 wire \mac2.sum_lvl2_ff[3] ;
 wire \mac2.sum_lvl2_ff[40] ;
 wire \mac2.sum_lvl2_ff[41] ;
 wire \mac2.sum_lvl2_ff[42] ;
 wire \mac2.sum_lvl2_ff[43] ;
 wire \mac2.sum_lvl2_ff[44] ;
 wire \mac2.sum_lvl2_ff[45] ;
 wire \mac2.sum_lvl2_ff[46] ;
 wire \mac2.sum_lvl2_ff[47] ;
 wire \mac2.sum_lvl2_ff[48] ;
 wire \mac2.sum_lvl2_ff[49] ;
 wire \mac2.sum_lvl2_ff[4] ;
 wire \mac2.sum_lvl2_ff[50] ;
 wire \mac2.sum_lvl2_ff[51] ;
 wire \mac2.sum_lvl2_ff[52] ;
 wire \mac2.sum_lvl2_ff[53] ;
 wire \mac2.sum_lvl2_ff[5] ;
 wire \mac2.sum_lvl2_ff[6] ;
 wire \mac2.sum_lvl2_ff[7] ;
 wire \mac2.sum_lvl2_ff[8] ;
 wire \mac2.sum_lvl2_ff[9] ;
 wire \mac2.sum_lvl3_ff[0] ;
 wire \mac2.sum_lvl3_ff[10] ;
 wire \mac2.sum_lvl3_ff[11] ;
 wire \mac2.sum_lvl3_ff[12] ;
 wire \mac2.sum_lvl3_ff[13] ;
 wire \mac2.sum_lvl3_ff[14] ;
 wire \mac2.sum_lvl3_ff[15] ;
 wire \mac2.sum_lvl3_ff[1] ;
 wire \mac2.sum_lvl3_ff[20] ;
 wire \mac2.sum_lvl3_ff[21] ;
 wire \mac2.sum_lvl3_ff[22] ;
 wire \mac2.sum_lvl3_ff[23] ;
 wire \mac2.sum_lvl3_ff[24] ;
 wire \mac2.sum_lvl3_ff[25] ;
 wire \mac2.sum_lvl3_ff[26] ;
 wire \mac2.sum_lvl3_ff[27] ;
 wire \mac2.sum_lvl3_ff[28] ;
 wire \mac2.sum_lvl3_ff[29] ;
 wire \mac2.sum_lvl3_ff[2] ;
 wire \mac2.sum_lvl3_ff[30] ;
 wire \mac2.sum_lvl3_ff[31] ;
 wire \mac2.sum_lvl3_ff[32] ;
 wire \mac2.sum_lvl3_ff[33] ;
 wire \mac2.sum_lvl3_ff[34] ;
 wire \mac2.sum_lvl3_ff[35] ;
 wire \mac2.sum_lvl3_ff[3] ;
 wire \mac2.sum_lvl3_ff[4] ;
 wire \mac2.sum_lvl3_ff[5] ;
 wire \mac2.sum_lvl3_ff[6] ;
 wire \mac2.sum_lvl3_ff[7] ;
 wire \mac2.sum_lvl3_ff[8] ;
 wire \mac2.sum_lvl3_ff[9] ;
 wire \mac2.total_sum[0] ;
 wire \mac2.total_sum[10] ;
 wire \mac2.total_sum[11] ;
 wire \mac2.total_sum[12] ;
 wire \mac2.total_sum[13] ;
 wire \mac2.total_sum[14] ;
 wire \mac2.total_sum[15] ;
 wire \mac2.total_sum[1] ;
 wire \mac2.total_sum[2] ;
 wire \mac2.total_sum[3] ;
 wire \mac2.total_sum[4] ;
 wire \mac2.total_sum[5] ;
 wire \mac2.total_sum[6] ;
 wire \mac2.total_sum[7] ;
 wire \mac2.total_sum[8] ;
 wire \mac2.total_sum[9] ;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_leaf_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net33;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;

 sg13g2_inv_1 _2983_ (.VDD(VPWR),
    .Y(_2587_),
    .A(\DP_3.I_range.out_data[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2984_ (.VDD(VPWR),
    .Y(_2588_),
    .A(\DP_3.I_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2985_ (.VDD(VPWR),
    .Y(_2589_),
    .A(\DP_3.Q_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2986_ (.VDD(VPWR),
    .Y(\DP_1.I_range.data_plus_4[6] ),
    .A(net4),
    .VSS(VGND));
 sg13g2_inv_1 _2987_ (.VDD(VPWR),
    .Y(\DP_3.I_range.data_plus_4[6] ),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _2988_ (.VDD(VPWR),
    .Y(\DP_3.Q_range.data_plus_4[6] ),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _2989_ (.VDD(VPWR),
    .Y(\DP_1.Q_range.data_plus_4[6] ),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _2990_ (.VDD(VPWR),
    .Y(_2590_),
    .A(net1010),
    .VSS(VGND));
 sg13g2_inv_1 _2991_ (.VDD(VPWR),
    .Y(_2591_),
    .A(net1005),
    .VSS(VGND));
 sg13g2_inv_1 _2992_ (.VDD(VPWR),
    .Y(_2592_),
    .A(net999),
    .VSS(VGND));
 sg13g2_inv_1 _2993_ (.VDD(VPWR),
    .Y(_2593_),
    .A(net995),
    .VSS(VGND));
 sg13g2_and2_1 _2994_ (.A(net958),
    .B(net903),
    .X(_0064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2995_ (.X(_2594_),
    .A(net956),
    .B(net898),
    .C(_0064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2996_ (.Y(_2595_),
    .B1(net898),
    .B2(net958),
    .A2(net956),
    .A1(net903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2997_ (.A(_2594_),
    .B(_2595_),
    .Y(_0065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2998_ (.A(net958),
    .B(net896),
    .X(_2596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2999_ (.A(net903),
    .B(net956),
    .C(net898),
    .D(net954),
    .X(_2597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3000_ (.Y(_2598_),
    .B1(net954),
    .B2(net903),
    .A2(net898),
    .A1(net956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3001_ (.A(_2597_),
    .B(_2598_),
    .Y(_2599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3002_ (.B(_2599_),
    .A(_2596_),
    .X(_2600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3003_ (.Y(_2601_),
    .A(_2594_),
    .B(_2600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3004_ (.B(_2600_),
    .A(_2594_),
    .X(_0066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3005_ (.Y(_2602_),
    .A(net958),
    .B(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2596_),
    .A2(_2599_),
    .Y(_2603_),
    .B1(_2597_));
 sg13g2_nand2_1 _3007_ (.Y(_2604_),
    .A(net956),
    .B(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3008_ (.A(net903),
    .B(net899),
    .C(net954),
    .D(net952),
    .X(_2605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3009_ (.B(net898),
    .C(net954),
    .A(net904),
    .Y(_2606_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net952));
 sg13g2_a22oi_1 _3010_ (.Y(_2607_),
    .B1(net952),
    .B2(net903),
    .A2(net954),
    .A1(net899),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3011_ (.A(_2604_),
    .B(_2605_),
    .C(_2607_),
    .Y(_2608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3012_ (.B1(_2604_),
    .VDD(VPWR),
    .Y(_2609_),
    .VSS(VGND),
    .A1(_2605_),
    .A2(_2607_));
 sg13g2_nor2b_1 _3013_ (.A(_2608_),
    .B_N(_2609_),
    .Y(_2610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3014_ (.Y(_2611_),
    .B(_2610_),
    .A_N(_2603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3015_ (.Y(_2612_),
    .A(_2603_),
    .B(_2610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3016_ (.Y(_2613_),
    .B(_2612_),
    .A_N(_2602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3017_ (.Y(_2614_),
    .A(_2602_),
    .B(_2612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3018_ (.A(_2601_),
    .B_N(_2614_),
    .Y(_2615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3019_ (.Y(_0067_),
    .A(_2601_),
    .B(_2614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3020_ (.Y(_2616_),
    .B1(net892),
    .B2(net958),
    .A2(net894),
    .A1(net956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3021_ (.Y(_2617_),
    .A(net956),
    .B(net892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3022_ (.A(_2602_),
    .B(_2617_),
    .Y(_2618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3023_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2619_),
    .B(_2618_),
    .A(_2616_));
 sg13g2_o21ai_1 _3024_ (.B1(_2606_),
    .VDD(VPWR),
    .Y(_2620_),
    .VSS(VGND),
    .A1(_2604_),
    .A2(_2607_));
 sg13g2_nand2_1 _3025_ (.Y(_2621_),
    .A(net954),
    .B(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3026_ (.A(net903),
    .B(net899),
    .C(net952),
    .D(net949),
    .X(_2622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3027_ (.B(net898),
    .C(net952),
    .A(net903),
    .Y(_2623_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net949));
 sg13g2_a22oi_1 _3028_ (.Y(_2624_),
    .B1(net949),
    .B2(net904),
    .A2(net952),
    .A1(net898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3029_ (.A(_2621_),
    .B(_2622_),
    .C(_2624_),
    .X(_2625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3030_ (.B1(_2621_),
    .VDD(VPWR),
    .Y(_2626_),
    .VSS(VGND),
    .A1(_2622_),
    .A2(_2624_));
 sg13g2_nand3_1 _3031_ (.B(_2625_),
    .C(_2626_),
    .A(_2620_),
    .Y(_2627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3032_ (.A2(_2626_),
    .A1(_2625_),
    .B1(_2620_),
    .X(_2628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3033_ (.Y(_2629_),
    .A(_2627_),
    .B(_2628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3034_ (.B(_2629_),
    .A(_2619_),
    .X(_2630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3035_ (.Y(_2631_),
    .A(_2611_),
    .B(_2613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3036_ (.Y(_2632_),
    .A(_2630_),
    .B(_2631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3037_ (.B(_2631_),
    .A(_2630_),
    .X(_2633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3038_ (.A(_2615_),
    .B(_2633_),
    .X(_2634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3039_ (.B(_2633_),
    .A(_2615_),
    .X(_0068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3040_ (.B1(_2627_),
    .VDD(VPWR),
    .Y(_2635_),
    .VSS(VGND),
    .A1(_2619_),
    .A2(_2629_));
 sg13g2_nand2_1 _3041_ (.Y(_2636_),
    .A(net958),
    .B(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3042_ (.Y(_2637_),
    .A(net955),
    .B(net892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3043_ (.Y(_2638_),
    .A(net954),
    .B(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3044_ (.B(_2638_),
    .A(_2617_),
    .X(_2639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3045_ (.Y(_2640_),
    .B(_2639_),
    .A_N(_2636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3046_ (.B(_2639_),
    .A(_2636_),
    .X(_2641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3047_ (.B1(_2623_),
    .VDD(VPWR),
    .Y(_2642_),
    .VSS(VGND),
    .A1(_2621_),
    .A2(_2624_));
 sg13g2_nand2_1 _3048_ (.Y(_2643_),
    .A(net896),
    .B(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3049_ (.A(net905),
    .B(net899),
    .C(net949),
    .D(net946),
    .X(_2644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3050_ (.B(net901),
    .C(net949),
    .A(net904),
    .Y(_2645_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net946));
 sg13g2_a22oi_1 _3051_ (.Y(_2646_),
    .B1(net946),
    .B2(net904),
    .A2(net949),
    .A1(net898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3052_ (.A(_2643_),
    .B(_2644_),
    .C(_2646_),
    .X(_2647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3053_ (.B1(_2643_),
    .VDD(VPWR),
    .Y(_2648_),
    .VSS(VGND),
    .A1(_2644_),
    .A2(_2646_));
 sg13g2_and3_1 _3054_ (.X(_2649_),
    .A(_2642_),
    .B(_2647_),
    .C(_2648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3055_ (.B(_2647_),
    .C(_2648_),
    .A(_2642_),
    .Y(_2650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3056_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2647_),
    .A2(_2648_),
    .Y(_2651_),
    .B1(_2642_));
 sg13g2_or3_1 _3057_ (.A(_2641_),
    .B(_2649_),
    .C(_2651_),
    .X(_2652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3058_ (.B1(_2641_),
    .VDD(VPWR),
    .Y(_2653_),
    .VSS(VGND),
    .A1(_2649_),
    .A2(_2651_));
 sg13g2_nand3_1 _3059_ (.B(_2652_),
    .C(_2653_),
    .A(_2635_),
    .Y(_2654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3060_ (.A2(_2653_),
    .A1(_2652_),
    .B1(_2635_),
    .X(_2655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3061_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2654_),
    .A2(_2655_),
    .Y(_2656_),
    .B1(_2618_));
 sg13g2_and3_1 _3062_ (.X(_2657_),
    .A(_2618_),
    .B(_2654_),
    .C(_2655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3063_ (.B(_2654_),
    .C(_2655_),
    .A(_2618_),
    .Y(_2658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3064_ (.A(_2632_),
    .B(_2656_),
    .C(_2657_),
    .Y(_2659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3065_ (.B1(_2632_),
    .VDD(VPWR),
    .Y(_2660_),
    .VSS(VGND),
    .A1(_2656_),
    .A2(_2657_));
 sg13g2_nand2b_1 _3066_ (.Y(_2661_),
    .B(_2660_),
    .A_N(_2659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3067_ (.Y(_0094_),
    .A(_2634_),
    .B(_2661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3068_ (.Y(_2662_),
    .A(_2654_),
    .B(_2658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3069_ (.B1(_2640_),
    .VDD(VPWR),
    .Y(_2663_),
    .VSS(VGND),
    .A1(_2617_),
    .A2(_2638_));
 sg13g2_nand2_2 _3070_ (.Y(_2664_),
    .A(net958),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3071_ (.Y(_2665_),
    .B(_2663_),
    .A_N(_2664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3072_ (.B(_2664_),
    .A(_2663_),
    .X(_2666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3073_ (.B1(_2650_),
    .VDD(VPWR),
    .Y(_2667_),
    .VSS(VGND),
    .A1(_2641_),
    .A2(_2651_));
 sg13g2_nand2_1 _3074_ (.Y(_2668_),
    .A(net956),
    .B(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3075_ (.Y(_2669_),
    .A(net953),
    .B(net892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3076_ (.Y(_2670_),
    .A(net952),
    .B(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3077_ (.B(_2670_),
    .A(_2637_),
    .X(_2671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3078_ (.Y(_2672_),
    .B(_2671_),
    .A_N(_2668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3079_ (.Y(_2673_),
    .A(_2668_),
    .B(_2671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3080_ (.B1(_2645_),
    .VDD(VPWR),
    .Y(_2674_),
    .VSS(VGND),
    .A1(_2643_),
    .A2(_2646_));
 sg13g2_nand2_1 _3081_ (.Y(_2675_),
    .A(net896),
    .B(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3082_ (.A(net904),
    .B(net901),
    .C(net946),
    .D(net944),
    .X(_2676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3083_ (.B(net900),
    .C(net946),
    .A(net904),
    .Y(_2677_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net944));
 sg13g2_a22oi_1 _3084_ (.Y(_2678_),
    .B1(net944),
    .B2(net904),
    .A2(net946),
    .A1(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3085_ (.A(_2675_),
    .B(_2676_),
    .C(_2678_),
    .X(_2679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3086_ (.B1(_2675_),
    .VDD(VPWR),
    .Y(_2680_),
    .VSS(VGND),
    .A1(_2676_),
    .A2(_2678_));
 sg13g2_and3_1 _3087_ (.X(_2681_),
    .A(_2674_),
    .B(_2679_),
    .C(_2680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3088_ (.B(_2679_),
    .C(_2680_),
    .A(_2674_),
    .Y(_2682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3089_ (.A2(_2680_),
    .A1(_2679_),
    .B1(_2674_),
    .X(_2683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3090_ (.B(_2682_),
    .C(_2683_),
    .A(_2673_),
    .Y(_2684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3091_ (.A2(_2683_),
    .A1(_2682_),
    .B1(_2673_),
    .X(_2685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3092_ (.B(_2684_),
    .C(_2685_),
    .A(_2667_),
    .Y(_2686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3093_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2684_),
    .A2(_2685_),
    .Y(_2687_),
    .B1(_2667_));
 sg13g2_a21o_1 _3094_ (.A2(_2685_),
    .A1(_2684_),
    .B1(_2667_),
    .X(_2688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3095_ (.Y(_2689_),
    .A(_2686_),
    .B(_2688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3096_ (.Y(_2690_),
    .A(_2666_),
    .B(_2689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3097_ (.Y(_2691_),
    .B(_2662_),
    .A_N(_2690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3098_ (.B(_2690_),
    .A(_2662_),
    .X(_2692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3099_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2634_),
    .A2(_2660_),
    .Y(_2693_),
    .B1(_2659_));
 sg13g2_xor2_1 _3100_ (.B(_2693_),
    .A(_2692_),
    .X(_0101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3101_ (.B1(_2686_),
    .VDD(VPWR),
    .Y(_2694_),
    .VSS(VGND),
    .A1(_2666_),
    .A2(_2687_));
 sg13g2_o21ai_1 _3102_ (.B1(_2672_),
    .VDD(VPWR),
    .Y(_2695_),
    .VSS(VGND),
    .A1(_2637_),
    .A2(_2670_));
 sg13g2_a22oi_1 _3103_ (.Y(_2696_),
    .B1(net887),
    .B2(net958),
    .A2(net889),
    .A1(net957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3104_ (.Y(_2697_),
    .A(net957),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3105_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2698_),
    .B(_2697_),
    .A(_2664_));
 sg13g2_nor2b_1 _3106_ (.A(_2696_),
    .B_N(_2698_),
    .Y(_2699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3107_ (.A(_2695_),
    .B(_2699_),
    .X(_2700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3108_ (.Y(_2701_),
    .A(_2695_),
    .B(_2699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3109_ (.A2(_2683_),
    .A1(_2673_),
    .B1(_2681_),
    .X(_2702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3110_ (.Y(_2703_),
    .A(net955),
    .B(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3111_ (.Y(_2704_),
    .A(net894),
    .B(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3112_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2705_),
    .B(_2704_),
    .A(_2669_));
 sg13g2_xnor2_1 _3113_ (.Y(_2706_),
    .A(_2669_),
    .B(_2704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3114_ (.Y(_2707_),
    .A(_2703_),
    .B(_2706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3115_ (.B1(_2677_),
    .VDD(VPWR),
    .Y(_2708_),
    .VSS(VGND),
    .A1(_2675_),
    .A2(_2678_));
 sg13g2_nand2_1 _3116_ (.Y(_2709_),
    .A(net896),
    .B(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3117_ (.A(net905),
    .B(net900),
    .C(net944),
    .D(net941),
    .X(_2710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3118_ (.B(net900),
    .C(net944),
    .A(net905),
    .Y(_2711_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net941));
 sg13g2_a22oi_1 _3119_ (.Y(_2712_),
    .B1(net941),
    .B2(net905),
    .A2(net944),
    .A1(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3120_ (.A(_2709_),
    .B(_2710_),
    .C(_2712_),
    .X(_2713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3121_ (.B1(_2709_),
    .VDD(VPWR),
    .Y(_2714_),
    .VSS(VGND),
    .A1(_2710_),
    .A2(_2712_));
 sg13g2_and3_1 _3122_ (.X(_2715_),
    .A(_2708_),
    .B(_2713_),
    .C(_2714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3123_ (.B(_2713_),
    .C(_2714_),
    .A(_2708_),
    .Y(_2716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3124_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2713_),
    .A2(_2714_),
    .Y(_2717_),
    .B1(_2708_));
 sg13g2_or3_1 _3125_ (.A(_2707_),
    .B(_2715_),
    .C(_2717_),
    .X(_2718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3126_ (.B1(_2707_),
    .VDD(VPWR),
    .Y(_2719_),
    .VSS(VGND),
    .A1(_2715_),
    .A2(_2717_));
 sg13g2_and3_1 _3127_ (.X(_2720_),
    .A(_2702_),
    .B(_2718_),
    .C(_2719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3128_ (.B(_2718_),
    .C(_2719_),
    .A(_2702_),
    .Y(_2721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3129_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2718_),
    .A2(_2719_),
    .Y(_2722_),
    .B1(_2702_));
 sg13g2_or3_1 _3130_ (.A(_2701_),
    .B(_2720_),
    .C(_2722_),
    .X(_2723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3131_ (.B1(_2701_),
    .VDD(VPWR),
    .Y(_2724_),
    .VSS(VGND),
    .A1(_2720_),
    .A2(_2722_));
 sg13g2_nand3_1 _3132_ (.B(_2723_),
    .C(_2724_),
    .A(_2694_),
    .Y(_2725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3133_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2723_),
    .A2(_2724_),
    .Y(_2726_),
    .B1(_2694_));
 sg13g2_a21o_1 _3134_ (.A2(_2724_),
    .A1(_2723_),
    .B1(_2694_),
    .X(_2727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3135_ (.Y(_2728_),
    .A(_2725_),
    .B(_2727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3136_ (.B(_2728_),
    .A(_2665_),
    .X(_2729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3137_ (.B1(_2691_),
    .VDD(VPWR),
    .Y(_2730_),
    .VSS(VGND),
    .A1(_2692_),
    .A2(_2693_));
 sg13g2_nand2_1 _3138_ (.Y(_2731_),
    .A(_2729_),
    .B(_2730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3139_ (.B(_2730_),
    .A(_2729_),
    .X(_0102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3140_ (.B1(_2721_),
    .VDD(VPWR),
    .Y(_2732_),
    .VSS(VGND),
    .A1(_2701_),
    .A2(_2722_));
 sg13g2_o21ai_1 _3141_ (.B1(_2705_),
    .VDD(VPWR),
    .Y(_2733_),
    .VSS(VGND),
    .A1(_2703_),
    .A2(_2706_));
 sg13g2_nand2_1 _3142_ (.Y(_2734_),
    .A(net959),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3143_ (.Y(_2735_),
    .A(net954),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3144_ (.Y(_2736_),
    .A(net955),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3145_ (.B(_2736_),
    .A(_2697_),
    .X(_2737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3146_ (.Y(_2738_),
    .B(_2737_),
    .A_N(_2734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3147_ (.Y(_2739_),
    .A(_2734_),
    .B(_2737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3148_ (.Y(_2740_),
    .A(_2733_),
    .B(_2739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3149_ (.Y(_2741_),
    .A(_2733_),
    .B(_2739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3150_ (.Y(_2742_),
    .A(_2698_),
    .B(_2741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3151_ (.B1(_2716_),
    .VDD(VPWR),
    .Y(_2743_),
    .VSS(VGND),
    .A1(_2707_),
    .A2(_2717_));
 sg13g2_nand2_1 _3152_ (.Y(_2744_),
    .A(net953),
    .B(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3153_ (.Y(_2745_),
    .A(net892),
    .B(net947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3154_ (.A(net894),
    .B(net950),
    .C(net892),
    .D(net946),
    .X(_2746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3155_ (.Y(_2747_),
    .B1(net947),
    .B2(net894),
    .A2(net892),
    .A1(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3156_ (.A(_2744_),
    .B(_2746_),
    .C(_2747_),
    .Y(_2748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3157_ (.B1(_2744_),
    .VDD(VPWR),
    .Y(_2749_),
    .VSS(VGND),
    .A1(_2746_),
    .A2(_2747_));
 sg13g2_nand2b_1 _3158_ (.Y(_2750_),
    .B(_2749_),
    .A_N(_2748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3159_ (.B1(_2711_),
    .VDD(VPWR),
    .Y(_2751_),
    .VSS(VGND),
    .A1(_2709_),
    .A2(_2712_));
 sg13g2_nand2_1 _3160_ (.Y(_2752_),
    .A(net896),
    .B(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3161_ (.A(net905),
    .B(net900),
    .C(net941),
    .D(net1006),
    .X(_2753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3162_ (.B(net900),
    .C(net941),
    .A(net905),
    .Y(_2754_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1006));
 sg13g2_a22oi_1 _3163_ (.Y(_2755_),
    .B1(net1006),
    .B2(net905),
    .A2(net941),
    .A1(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3164_ (.A(_2752_),
    .B(_2753_),
    .C(_2755_),
    .X(_2756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3165_ (.B1(_2752_),
    .VDD(VPWR),
    .Y(_2757_),
    .VSS(VGND),
    .A1(_2753_),
    .A2(_2755_));
 sg13g2_and3_1 _3166_ (.X(_2758_),
    .A(_2751_),
    .B(_2756_),
    .C(_2757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3167_ (.B(_2756_),
    .C(_2757_),
    .A(_2751_),
    .Y(_2759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2756_),
    .A2(_2757_),
    .Y(_2760_),
    .B1(_2751_));
 sg13g2_or3_1 _3169_ (.A(_2750_),
    .B(_2758_),
    .C(_2760_),
    .X(_2761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3170_ (.B1(_2750_),
    .VDD(VPWR),
    .Y(_2762_),
    .VSS(VGND),
    .A1(_2758_),
    .A2(_2760_));
 sg13g2_and3_1 _3171_ (.X(_2763_),
    .A(_2743_),
    .B(_2761_),
    .C(_2762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3172_ (.B(_2761_),
    .C(_2762_),
    .A(_2743_),
    .Y(_2764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3173_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2761_),
    .A2(_2762_),
    .Y(_2765_),
    .B1(_2743_));
 sg13g2_or3_1 _3174_ (.A(_2742_),
    .B(_2763_),
    .C(_2765_),
    .X(_2766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3175_ (.B1(_2742_),
    .VDD(VPWR),
    .Y(_2767_),
    .VSS(VGND),
    .A1(_2763_),
    .A2(_2765_));
 sg13g2_nand3_1 _3176_ (.B(_2766_),
    .C(_2767_),
    .A(_2732_),
    .Y(_2768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3177_ (.A2(_2767_),
    .A1(_2766_),
    .B1(_2732_),
    .X(_2769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3178_ (.A2(_2769_),
    .A1(_2768_),
    .B1(_2700_),
    .X(_2770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3179_ (.B(_2768_),
    .C(_2769_),
    .A(_2700_),
    .Y(_2771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3180_ (.B1(_2725_),
    .VDD(VPWR),
    .Y(_2772_),
    .VSS(VGND),
    .A1(_2665_),
    .A2(_2726_));
 sg13g2_nand3_1 _3181_ (.B(_2771_),
    .C(_2772_),
    .A(_2770_),
    .Y(_2773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3182_ (.A2(_2771_),
    .A1(_2770_),
    .B1(_2772_),
    .X(_2774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3183_ (.A(_2773_),
    .B(_2774_),
    .X(_2775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3184_ (.B(_2730_),
    .C(_2775_),
    .A(_2729_),
    .Y(_2776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3185_ (.Y(_0103_),
    .A(_2731_),
    .B(_2775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3186_ (.B1(_2740_),
    .VDD(VPWR),
    .Y(_2777_),
    .VSS(VGND),
    .A1(_2698_),
    .A2(_2741_));
 sg13g2_o21ai_1 _3187_ (.B1(_2764_),
    .VDD(VPWR),
    .Y(_2778_),
    .VSS(VGND),
    .A1(_2742_),
    .A2(_2765_));
 sg13g2_o21ai_1 _3188_ (.B1(_2738_),
    .VDD(VPWR),
    .Y(_2779_),
    .VSS(VGND),
    .A1(_2697_),
    .A2(_2736_));
 sg13g2_or2_1 _3189_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2780_),
    .B(_2748_),
    .A(_2746_));
 sg13g2_nand2_1 _3190_ (.Y(_2781_),
    .A(net957),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3191_ (.Y(_2782_),
    .A(net953),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3192_ (.Y(_2783_),
    .A(net953),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3193_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2784_),
    .B(_2782_),
    .A(_2736_));
 sg13g2_xnor2_1 _3194_ (.Y(_2785_),
    .A(_2735_),
    .B(_2783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3195_ (.B(_2785_),
    .A(_2781_),
    .X(_2786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3196_ (.Y(_2787_),
    .A(_2780_),
    .B(_2786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3197_ (.A(_2787_),
    .B_N(_2779_),
    .Y(_2788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3198_ (.B(_2787_),
    .A(_2779_),
    .X(_2789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3199_ (.B1(_2759_),
    .VDD(VPWR),
    .Y(_2790_),
    .VSS(VGND),
    .A1(_2750_),
    .A2(_2760_));
 sg13g2_nand2_1 _3200_ (.Y(_2791_),
    .A(net950),
    .B(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3201_ (.Y(_2792_),
    .A(net894),
    .B(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3202_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2793_),
    .B(_2792_),
    .A(_2745_));
 sg13g2_and2_1 _3203_ (.A(_2745_),
    .B(_2792_),
    .X(_2794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3204_ (.Y(_2795_),
    .A(_2745_),
    .B(_2792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3205_ (.Y(_2796_),
    .A(_2791_),
    .B(_2795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3206_ (.B1(_2754_),
    .VDD(VPWR),
    .Y(_2797_),
    .VSS(VGND),
    .A1(_2752_),
    .A2(_2755_));
 sg13g2_nand2_1 _3207_ (.Y(_2798_),
    .A(net896),
    .B(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3208_ (.A(net901),
    .B(net897),
    .C(net941),
    .D(net1006),
    .X(_2799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3209_ (.Y(_2800_),
    .B1(net1006),
    .B2(net901),
    .A2(net942),
    .A1(net897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3210_ (.A(_2799_),
    .B(_2800_),
    .Y(_2801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3211_ (.Y(_2802_),
    .A(_2797_),
    .B(_2801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3212_ (.Y(_2803_),
    .A(_2797_),
    .B(_2801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3213_ (.B(_2803_),
    .A(_2796_),
    .X(_2804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3214_ (.Y(_2805_),
    .A(_2790_),
    .B(_2804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3215_ (.Y(_2806_),
    .A(_2790_),
    .B(_2804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3216_ (.B(_2806_),
    .A(_2789_),
    .X(_2807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3217_ (.Y(_2808_),
    .A(_2778_),
    .B(_2807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3218_ (.Y(_2809_),
    .A(_2778_),
    .B(_2807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3219_ (.Y(_2810_),
    .B(_2777_),
    .A_N(_2809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3220_ (.B(_2809_),
    .A(_2777_),
    .X(_2811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3221_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2768_),
    .A2(_2771_),
    .Y(_2812_),
    .B1(_2811_));
 sg13g2_a21o_1 _3222_ (.A2(_2771_),
    .A1(_2768_),
    .B1(_2811_),
    .X(_2813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3223_ (.X(_2814_),
    .A(_2768_),
    .B(_2771_),
    .C(_2811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3224_ (.A(_2812_),
    .B(_2814_),
    .Y(_2815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3225_ (.Y(_2816_),
    .A(_2773_),
    .B(_2776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3226_ (.B(_2816_),
    .A(_2815_),
    .X(_0104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3227_ (.A2(_2786_),
    .A1(_2780_),
    .B1(_2788_),
    .X(_2817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3228_ (.B1(_2805_),
    .VDD(VPWR),
    .Y(_2818_),
    .VSS(VGND),
    .A1(_2789_),
    .A2(_2806_));
 sg13g2_o21ai_1 _3229_ (.B1(_2784_),
    .VDD(VPWR),
    .Y(_2819_),
    .VSS(VGND),
    .A1(_2781_),
    .A2(_2785_));
 sg13g2_o21ai_1 _3230_ (.B1(_2793_),
    .VDD(VPWR),
    .Y(_2820_),
    .VSS(VGND),
    .A1(_2791_),
    .A2(_2794_));
 sg13g2_nand2_1 _3231_ (.Y(_2821_),
    .A(net955),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3232_ (.Y(_2822_),
    .A(net949),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3233_ (.Y(_2823_),
    .A(net950),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3234_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2824_),
    .B(_2822_),
    .A(_2783_));
 sg13g2_xnor2_1 _3235_ (.Y(_2825_),
    .A(_2782_),
    .B(_2823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3236_ (.B(_2825_),
    .A(_2821_),
    .X(_2826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3237_ (.Y(_2827_),
    .A(_2820_),
    .B(_2826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3238_ (.A(_2827_),
    .B_N(_2819_),
    .Y(_2828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3239_ (.B(_2827_),
    .A(_2819_),
    .X(_2829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3240_ (.B1(_2802_),
    .VDD(VPWR),
    .Y(_2830_),
    .VSS(VGND),
    .A1(_2796_),
    .A2(_2803_));
 sg13g2_a21oi_1 _3241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net901),
    .A2(net942),
    .Y(_2831_),
    .B1(_2798_));
 sg13g2_nand2_1 _3242_ (.Y(_2832_),
    .A(net947),
    .B(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3243_ (.Y(_2833_),
    .A(net893),
    .B(net943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3244_ (.A(net895),
    .B(net892),
    .C(net945),
    .D(net942),
    .X(_2834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3245_ (.Y(_2835_),
    .B1(net941),
    .B2(net895),
    .A2(net945),
    .A1(net893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3246_ (.A(_2832_),
    .B(_2834_),
    .C(_2835_),
    .Y(_2836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3247_ (.B1(_2832_),
    .VDD(VPWR),
    .Y(_2837_),
    .VSS(VGND),
    .A1(_2834_),
    .A2(_2835_));
 sg13g2_nor2b_1 _3248_ (.A(_2836_),
    .B_N(_2837_),
    .Y(_2838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3249_ (.Y(_2839_),
    .A(_2831_),
    .B(_2838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3250_ (.Y(_2840_),
    .B(_2830_),
    .A_N(_2839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3251_ (.B(_2839_),
    .A(_2830_),
    .X(_2841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3252_ (.B(_2841_),
    .A(_2829_),
    .X(_2842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3253_ (.Y(_2843_),
    .A(_2818_),
    .B(_2842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3254_ (.B(_2842_),
    .A(_2818_),
    .X(_2844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3255_ (.Y(_2845_),
    .A(_2817_),
    .B(_2844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3256_ (.Y(_2846_),
    .A(_2817_),
    .B(_2844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3257_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2808_),
    .A2(_2810_),
    .Y(_2847_),
    .B1(_2846_));
 sg13g2_nand3_1 _3258_ (.B(_2810_),
    .C(_2846_),
    .A(_2808_),
    .Y(_2848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3259_ (.A(_2847_),
    .B_N(_2848_),
    .Y(_2849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3260_ (.B(_2730_),
    .C(_2775_),
    .A(_2729_),
    .Y(_2850_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2815_));
 sg13g2_a21oi_1 _3261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2773_),
    .A2(_2813_),
    .Y(_2851_),
    .B1(_2814_));
 sg13g2_nand2b_1 _3262_ (.Y(_2852_),
    .B(_2850_),
    .A_N(_2851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3263_ (.B(_2852_),
    .A(_2849_),
    .X(_0095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3264_ (.A2(_2826_),
    .A1(_2820_),
    .B1(_2828_),
    .X(_2853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3265_ (.B1(_2840_),
    .VDD(VPWR),
    .Y(_2854_),
    .VSS(VGND),
    .A1(_2829_),
    .A2(_2841_));
 sg13g2_a21o_1 _3266_ (.A2(_2838_),
    .A1(_2831_),
    .B1(_2799_),
    .X(_2855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3267_ (.Y(_2856_),
    .A(net890),
    .B(net945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3268_ (.Y(_2857_),
    .A(net895),
    .B(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3269_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2858_),
    .B(_2857_),
    .A(_2833_));
 sg13g2_xnor2_1 _3270_ (.Y(_2859_),
    .A(_2833_),
    .B(_2857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3271_ (.B(_2859_),
    .A(_2856_),
    .X(_2860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3272_ (.Y(_2861_),
    .A(_2855_),
    .B(_2860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3273_ (.B1(_2824_),
    .VDD(VPWR),
    .Y(_2862_),
    .VSS(VGND),
    .A1(_2821_),
    .A2(_2825_));
 sg13g2_or2_1 _3274_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2863_),
    .B(_2836_),
    .A(_2834_));
 sg13g2_nand2_1 _3275_ (.Y(_2864_),
    .A(net953),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3276_ (.Y(_2865_),
    .A(net948),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3277_ (.Y(_2866_),
    .A(net947),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3278_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2867_),
    .B(_2865_),
    .A(_2823_));
 sg13g2_xnor2_1 _3279_ (.Y(_2868_),
    .A(_2822_),
    .B(_2866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3280_ (.B(_2868_),
    .A(_2864_),
    .X(_2869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3281_ (.Y(_2870_),
    .A(_2863_),
    .B(_2869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3282_ (.A(_2870_),
    .B_N(_2862_),
    .Y(_2871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3283_ (.B(_2870_),
    .A(_2862_),
    .X(_2872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3284_ (.A(_2861_),
    .B(_2872_),
    .Y(_2873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3285_ (.B(_2872_),
    .A(_2861_),
    .X(_2874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3286_ (.Y(_2875_),
    .A(_2854_),
    .B(_2874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3287_ (.A(_2875_),
    .B_N(_2853_),
    .Y(_2876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3288_ (.B(_2875_),
    .A(_2853_),
    .X(_2877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3289_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2843_),
    .A2(_2845_),
    .Y(_2878_),
    .B1(_2877_));
 sg13g2_nand3_1 _3290_ (.B(_2845_),
    .C(_2877_),
    .A(_2843_),
    .Y(_2879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3291_ (.A(_2878_),
    .B_N(_2879_),
    .Y(_2880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3292_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2849_),
    .A2(_2852_),
    .Y(_2881_),
    .B1(_2847_));
 sg13g2_xnor2_1 _3293_ (.Y(_0096_),
    .A(_2880_),
    .B(_2881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3294_ (.A2(_2869_),
    .A1(_2863_),
    .B1(_2871_),
    .X(_2882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3295_ (.Y(_2883_),
    .B1(net1007),
    .B2(net893),
    .A2(net943),
    .A1(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3296_ (.Y(_2884_),
    .A(net891),
    .B(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3297_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2885_),
    .B(_2884_),
    .A(_2833_));
 sg13g2_nand2b_1 _3298_ (.Y(_2886_),
    .B(_2885_),
    .A_N(_2883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3299_ (.B1(_2867_),
    .VDD(VPWR),
    .Y(_2887_),
    .VSS(VGND),
    .A1(_2864_),
    .A2(_2868_));
 sg13g2_o21ai_1 _3300_ (.B1(_2858_),
    .VDD(VPWR),
    .Y(_2888_),
    .VSS(VGND),
    .A1(_2856_),
    .A2(_2859_));
 sg13g2_nand2_1 _3301_ (.Y(_2889_),
    .A(net951),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3302_ (.Y(_2890_),
    .A(net945),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3303_ (.Y(_2891_),
    .A(net945),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3304_ (.B(_2891_),
    .A(_2865_),
    .X(_2892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3305_ (.Y(_2893_),
    .B(_2892_),
    .A_N(_2889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3306_ (.Y(_2894_),
    .A(_2889_),
    .B(_2892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3307_ (.Y(_2895_),
    .A(_2888_),
    .B(_2894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3308_ (.A(_2895_),
    .B_N(_2887_),
    .Y(_2896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3309_ (.B(_2895_),
    .A(_2887_),
    .X(_2897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3310_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2898_),
    .B(_2897_),
    .A(_2886_));
 sg13g2_xor2_1 _3311_ (.B(_2897_),
    .A(_2886_),
    .X(_2899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3312_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2855_),
    .A2(_2860_),
    .Y(_2900_),
    .B1(_2873_));
 sg13g2_nor2b_1 _3313_ (.A(_2900_),
    .B_N(_2899_),
    .Y(_2901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3314_ (.Y(_2902_),
    .A(_2899_),
    .B(_2900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3315_ (.Y(_2903_),
    .A(_2882_),
    .B(_2902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3316_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2854_),
    .A2(_2874_),
    .Y(_2904_),
    .B1(_2876_));
 sg13g2_or2_1 _3317_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2905_),
    .B(_2904_),
    .A(_2903_));
 sg13g2_xor2_1 _3318_ (.B(_2904_),
    .A(_2903_),
    .X(_2906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3319_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2847_),
    .A2(_2879_),
    .Y(_2907_),
    .B1(_2878_));
 sg13g2_nor2b_1 _3320_ (.A(_2851_),
    .B_N(_2907_),
    .Y(_2908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3321_ (.B1(_2879_),
    .VDD(VPWR),
    .Y(_2909_),
    .VSS(VGND),
    .A1(_2848_),
    .A2(_2878_));
 sg13g2_a21oi_2 _3322_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2909_),
    .Y(_2910_),
    .A2(_2908_),
    .A1(_2850_));
 sg13g2_nand2_1 _3323_ (.Y(_2911_),
    .A(_2906_),
    .B(_2910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3324_ (.B(_2910_),
    .A(_2906_),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3325_ (.A2(_2902_),
    .A1(_2882_),
    .B1(_2901_),
    .X(_2912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3326_ (.A2(_2894_),
    .A1(_2888_),
    .B1(_2896_),
    .X(_2913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3327_ (.B1(_2893_),
    .VDD(VPWR),
    .Y(_2914_),
    .VSS(VGND),
    .A1(_2865_),
    .A2(_2891_));
 sg13g2_nand2_1 _3328_ (.Y(_2915_),
    .A(net948),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3329_ (.Y(_2916_),
    .A(net943),
    .B(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3330_ (.Y(_2917_),
    .A(net889),
    .B(net943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3331_ (.B(_2917_),
    .A(_2890_),
    .X(_2918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3332_ (.Y(_2919_),
    .B(_2918_),
    .A_N(_2915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3333_ (.Y(_2920_),
    .A(_2915_),
    .B(_2918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3334_ (.A(_2885_),
    .B_N(_2920_),
    .Y(_2921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3335_ (.Y(_2922_),
    .A(_2885_),
    .B(_2920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3336_ (.Y(_2923_),
    .A(_2914_),
    .B(_2922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3337_ (.A(_2884_),
    .B(_2923_),
    .Y(_2924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3338_ (.B(_2923_),
    .A(_2884_),
    .X(_2925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3339_ (.Y(_2926_),
    .B(_2925_),
    .A_N(_2898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3340_ (.Y(_2927_),
    .A(_2898_),
    .B(_2925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3341_ (.Y(_2928_),
    .A(_2913_),
    .B(_2927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3342_ (.B(_2927_),
    .A(_2913_),
    .X(_2929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3343_ (.Y(_2930_),
    .A(_2912_),
    .B(_2929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3344_ (.A(_2912_),
    .B(_2929_),
    .Y(_2931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3345_ (.B(_2929_),
    .A(_2912_),
    .X(_2932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3346_ (.Y(_2933_),
    .A(_2905_),
    .B(_2911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3347_ (.B(_2933_),
    .A(_2932_),
    .X(_0098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3348_ (.A(_2906_),
    .B(_2932_),
    .X(_2934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3349_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2905_),
    .A2(_2930_),
    .Y(_2935_),
    .B1(_2931_));
 sg13g2_a21o_1 _3350_ (.A2(_2934_),
    .A1(_2910_),
    .B1(_2935_),
    .X(_2936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3351_ (.A(_2926_),
    .B(_2928_),
    .X(_2937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3352_ (.A2(_2922_),
    .A1(_2914_),
    .B1(_2921_),
    .X(_2938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3353_ (.Y(_2939_),
    .A(net945),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3354_ (.Y(_2940_),
    .A(net888),
    .B(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3355_ (.Y(_2941_),
    .A(\DP_2.matrix[78] ),
    .B(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3356_ (.B(_2941_),
    .A(_2916_),
    .X(_2942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3357_ (.Y(_2943_),
    .B(_2942_),
    .A_N(_2939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3358_ (.Y(_2944_),
    .A(_2939_),
    .B(_2942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3359_ (.B1(_2919_),
    .VDD(VPWR),
    .Y(_2945_),
    .VSS(VGND),
    .A1(_2890_),
    .A2(_2917_));
 sg13g2_nand2_1 _3360_ (.Y(_2946_),
    .A(_2944_),
    .B(_2945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3361_ (.B(_2945_),
    .A(_2944_),
    .X(_2947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3362_ (.Y(_2948_),
    .A(_2924_),
    .B(_2947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3363_ (.A(_2948_),
    .B_N(_2938_),
    .Y(_2949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3364_ (.B(_2948_),
    .A(_2938_),
    .X(_2950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3365_ (.A(_2937_),
    .B(_2950_),
    .Y(_2951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3366_ (.B(_2950_),
    .A(_2937_),
    .X(_2952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3367_ (.B(_2952_),
    .A(_2936_),
    .X(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3368_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2936_),
    .A2(_2952_),
    .Y(_2953_),
    .B1(_2951_));
 sg13g2_a21oi_1 _3369_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2924_),
    .A2(_2947_),
    .Y(_2954_),
    .B1(_2949_));
 sg13g2_o21ai_1 _3370_ (.B1(_2943_),
    .VDD(VPWR),
    .Y(_2955_),
    .VSS(VGND),
    .A1(_2917_),
    .A2(_2940_));
 sg13g2_nand2_1 _3371_ (.Y(_2956_),
    .A(net943),
    .B(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3372_ (.Y(_2957_),
    .A(_2940_),
    .B(_2956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3373_ (.Y(_2958_),
    .A(_2955_),
    .B(_2957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3374_ (.Y(_2959_),
    .A(_2946_),
    .B(_2958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3375_ (.Y(_2960_),
    .A(_2954_),
    .B(_2959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3376_ (.Y(_0100_),
    .A(_2953_),
    .B(_2960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3377_ (.A(net993),
    .B(net937),
    .X(_0069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3378_ (.X(_2961_),
    .A(net991),
    .B(net932),
    .C(_0069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3379_ (.Y(_2962_),
    .B1(net932),
    .B2(net993),
    .A2(net991),
    .A1(net937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3380_ (.A(_2961_),
    .B(_2962_),
    .Y(_0070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3381_ (.A(net993),
    .B(net930),
    .X(_2963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3382_ (.A(net937),
    .B(net991),
    .C(net932),
    .D(net989),
    .X(_2964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3383_ (.Y(_2965_),
    .B1(net989),
    .B2(net940),
    .A2(net936),
    .A1(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3384_ (.A(_2964_),
    .B(_2965_),
    .Y(_2966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3385_ (.B(_2966_),
    .A(_2963_),
    .X(_2967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3386_ (.Y(_2968_),
    .A(_2961_),
    .B(_2967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3387_ (.B(_2967_),
    .A(_2961_),
    .X(_0071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3388_ (.Y(_2969_),
    .A(net358),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3389_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2963_),
    .A2(_2966_),
    .Y(_2970_),
    .B1(_2964_));
 sg13g2_nand2_1 _3390_ (.Y(_2971_),
    .A(net991),
    .B(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3391_ (.A(net937),
    .B(net932),
    .C(net989),
    .D(net987),
    .X(_2972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3392_ (.B(net932),
    .C(net989),
    .A(net940),
    .Y(_2973_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net987));
 sg13g2_a22oi_1 _3393_ (.Y(_2974_),
    .B1(net987),
    .B2(net937),
    .A2(net989),
    .A1(net932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3394_ (.A(_2971_),
    .B(_2972_),
    .C(_2974_),
    .Y(_2975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3395_ (.B1(_2971_),
    .VDD(VPWR),
    .Y(_2976_),
    .VSS(VGND),
    .A1(_2972_),
    .A2(_2974_));
 sg13g2_nor2b_1 _3396_ (.A(_2975_),
    .B_N(_2976_),
    .Y(_2977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3397_ (.Y(_2978_),
    .B(_2977_),
    .A_N(_2970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3398_ (.Y(_2979_),
    .A(_2970_),
    .B(_2977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3399_ (.Y(_2980_),
    .B(_2979_),
    .A_N(_2969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3400_ (.Y(_2981_),
    .A(_2969_),
    .B(_2979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3401_ (.A(_2968_),
    .B_N(_2981_),
    .Y(_2982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3402_ (.Y(_0072_),
    .A(_2968_),
    .B(_2981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3403_ (.Y(_0268_),
    .B1(net928),
    .B2(net993),
    .A2(net929),
    .A1(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3404_ (.Y(_0269_),
    .A(net992),
    .B(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3405_ (.A(_2969_),
    .B(_0269_),
    .Y(_0270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3406_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0271_),
    .B(_0270_),
    .A(_0268_));
 sg13g2_o21ai_1 _3407_ (.B1(_2973_),
    .VDD(VPWR),
    .Y(_0272_),
    .VSS(VGND),
    .A1(_2971_),
    .A2(_2974_));
 sg13g2_nand2_1 _3408_ (.Y(_0273_),
    .A(net989),
    .B(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3409_ (.A(net937),
    .B(net936),
    .C(net987),
    .D(net985),
    .X(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3410_ (.B(net935),
    .C(net987),
    .A(net939),
    .Y(_0275_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net985));
 sg13g2_a22oi_1 _3411_ (.Y(_0276_),
    .B1(net985),
    .B2(net939),
    .A2(net987),
    .A1(net936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3412_ (.A(_0273_),
    .B(_0274_),
    .C(_0276_),
    .X(_0277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3413_ (.B1(_0273_),
    .VDD(VPWR),
    .Y(_0278_),
    .VSS(VGND),
    .A1(_0274_),
    .A2(_0276_));
 sg13g2_nand3_1 _3414_ (.B(_0277_),
    .C(_0278_),
    .A(_0272_),
    .Y(_0279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3415_ (.A2(_0278_),
    .A1(_0277_),
    .B1(_0272_),
    .X(_0280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3416_ (.Y(_0281_),
    .A(_0279_),
    .B(_0280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3417_ (.B(_0281_),
    .A(_0271_),
    .X(_0282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3418_ (.Y(_0283_),
    .A(_2978_),
    .B(_2980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3419_ (.Y(_0284_),
    .A(_0282_),
    .B(_0283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3420_ (.B(_0283_),
    .A(_0282_),
    .X(_0285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3421_ (.A(_2982_),
    .B(_0285_),
    .X(_0286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3422_ (.B(_0285_),
    .A(_2982_),
    .X(_0073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3423_ (.B1(_0279_),
    .VDD(VPWR),
    .Y(_0287_),
    .VSS(VGND),
    .A1(_0271_),
    .A2(_0281_));
 sg13g2_nand2_1 _3424_ (.Y(_0288_),
    .A(net993),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3425_ (.Y(_0289_),
    .A(net990),
    .B(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3426_ (.Y(_0290_),
    .A(net990),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3427_ (.B(_0290_),
    .A(_0269_),
    .X(_0291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3428_ (.Y(_0292_),
    .B(_0291_),
    .A_N(_0288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3429_ (.B(_0291_),
    .A(_0288_),
    .X(_0293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3430_ (.B1(_0275_),
    .VDD(VPWR),
    .Y(_0294_),
    .VSS(VGND),
    .A1(_0273_),
    .A2(_0276_));
 sg13g2_nand2_1 _3431_ (.Y(_0295_),
    .A(net931),
    .B(net988),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3432_ (.A(net939),
    .B(net935),
    .C(net985),
    .D(net983),
    .X(_0296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3433_ (.B(net935),
    .C(net985),
    .A(net939),
    .Y(_0297_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net983));
 sg13g2_a22oi_1 _3434_ (.Y(_0298_),
    .B1(net983),
    .B2(net939),
    .A2(net985),
    .A1(net935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3435_ (.A(_0295_),
    .B(_0296_),
    .C(_0298_),
    .X(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3436_ (.B1(_0295_),
    .VDD(VPWR),
    .Y(_0300_),
    .VSS(VGND),
    .A1(_0296_),
    .A2(_0298_));
 sg13g2_and3_1 _3437_ (.X(_0301_),
    .A(_0294_),
    .B(_0299_),
    .C(_0300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3438_ (.B(_0299_),
    .C(_0300_),
    .A(_0294_),
    .Y(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0299_),
    .A2(_0300_),
    .Y(_0303_),
    .B1(_0294_));
 sg13g2_or3_1 _3440_ (.A(_0293_),
    .B(_0301_),
    .C(_0303_),
    .X(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3441_ (.B1(_0293_),
    .VDD(VPWR),
    .Y(_0305_),
    .VSS(VGND),
    .A1(_0301_),
    .A2(_0303_));
 sg13g2_nand3_1 _3442_ (.B(_0304_),
    .C(_0305_),
    .A(_0287_),
    .Y(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3443_ (.A2(_0305_),
    .A1(_0304_),
    .B1(_0287_),
    .X(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3444_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0306_),
    .A2(_0307_),
    .Y(_0308_),
    .B1(_0270_));
 sg13g2_and3_1 _3445_ (.X(_0309_),
    .A(_0270_),
    .B(_0306_),
    .C(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3446_ (.B(_0306_),
    .C(_0307_),
    .A(_0270_),
    .Y(_0310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3447_ (.A(_0284_),
    .B(_0308_),
    .C(_0309_),
    .Y(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3448_ (.B1(_0284_),
    .VDD(VPWR),
    .Y(_0312_),
    .VSS(VGND),
    .A1(_0308_),
    .A2(_0309_));
 sg13g2_nand2b_1 _3449_ (.Y(_0313_),
    .B(_0312_),
    .A_N(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3450_ (.Y(_0105_),
    .A(_0286_),
    .B(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3451_ (.Y(_0314_),
    .A(_0306_),
    .B(_0310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3452_ (.B1(_0292_),
    .VDD(VPWR),
    .Y(_0315_),
    .VSS(VGND),
    .A1(_0269_),
    .A2(_0290_));
 sg13g2_nand2_1 _3453_ (.Y(_0316_),
    .A(\DP_1.matrix[0] ),
    .B(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3454_ (.Y(_0317_),
    .B(_0315_),
    .A_N(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3455_ (.B(_0316_),
    .A(_0315_),
    .X(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3456_ (.B1(_0302_),
    .VDD(VPWR),
    .Y(_0319_),
    .VSS(VGND),
    .A1(_0293_),
    .A2(_0303_));
 sg13g2_nand2_1 _3457_ (.Y(_0320_),
    .A(net991),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3458_ (.Y(_0321_),
    .A(net988),
    .B(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3459_ (.Y(_0322_),
    .A(net988),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3460_ (.B(_0322_),
    .A(_0289_),
    .X(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3461_ (.Y(_0324_),
    .B(_0323_),
    .A_N(_0320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3462_ (.Y(_0325_),
    .A(_0320_),
    .B(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3463_ (.B1(_0297_),
    .VDD(VPWR),
    .Y(_0326_),
    .VSS(VGND),
    .A1(_0295_),
    .A2(_0298_));
 sg13g2_nand2_1 _3464_ (.Y(_0327_),
    .A(net931),
    .B(net986),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3465_ (.A(net938),
    .B(net935),
    .C(net983),
    .D(net981),
    .X(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3466_ (.B(net933),
    .C(net983),
    .A(net938),
    .Y(_0329_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net981));
 sg13g2_a22oi_1 _3467_ (.Y(_0330_),
    .B1(net981),
    .B2(net938),
    .A2(net983),
    .A1(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3468_ (.A(_0327_),
    .B(_0328_),
    .C(_0330_),
    .X(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3469_ (.B1(_0327_),
    .VDD(VPWR),
    .Y(_0332_),
    .VSS(VGND),
    .A1(_0328_),
    .A2(_0330_));
 sg13g2_and3_1 _3470_ (.X(_0333_),
    .A(_0326_),
    .B(_0331_),
    .C(_0332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3471_ (.B(_0331_),
    .C(_0332_),
    .A(_0326_),
    .Y(_0334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3472_ (.A2(_0332_),
    .A1(_0331_),
    .B1(_0326_),
    .X(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3473_ (.B(_0334_),
    .C(_0335_),
    .A(_0325_),
    .Y(_0336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3474_ (.A2(_0335_),
    .A1(_0334_),
    .B1(_0325_),
    .X(_0337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3475_ (.B(_0336_),
    .C(_0337_),
    .A(_0319_),
    .Y(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3476_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0336_),
    .A2(_0337_),
    .Y(_0339_),
    .B1(_0319_));
 sg13g2_a21o_1 _3477_ (.A2(_0337_),
    .A1(_0336_),
    .B1(_0319_),
    .X(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3478_ (.Y(_0341_),
    .A(_0338_),
    .B(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3479_ (.Y(_0342_),
    .A(_0318_),
    .B(_0341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3480_ (.Y(_0343_),
    .B(_0314_),
    .A_N(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3481_ (.B(_0342_),
    .A(_0314_),
    .X(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3482_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0286_),
    .A2(_0312_),
    .Y(_0345_),
    .B1(_0311_));
 sg13g2_xor2_1 _3483_ (.B(_0345_),
    .A(_0344_),
    .X(_0112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3484_ (.B1(_0338_),
    .VDD(VPWR),
    .Y(_0346_),
    .VSS(VGND),
    .A1(_0318_),
    .A2(_0339_));
 sg13g2_o21ai_1 _3485_ (.B1(_0324_),
    .VDD(VPWR),
    .Y(_0347_),
    .VSS(VGND),
    .A1(_0289_),
    .A2(_0322_));
 sg13g2_a22oi_1 _3486_ (.Y(_0348_),
    .B1(net925),
    .B2(net993),
    .A2(net926),
    .A1(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3487_ (.Y(_0349_),
    .A(net992),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3488_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0350_),
    .B(_0349_),
    .A(_0316_));
 sg13g2_nor2b_1 _3489_ (.A(_0348_),
    .B_N(_0350_),
    .Y(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3490_ (.A(_0347_),
    .B(_0351_),
    .X(_0352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3491_ (.Y(_0353_),
    .A(_0347_),
    .B(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3492_ (.A2(_0335_),
    .A1(_0325_),
    .B1(_0333_),
    .X(_0354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3493_ (.Y(_0355_),
    .A(net990),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3494_ (.Y(_0356_),
    .A(net986),
    .B(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3495_ (.Y(_0357_),
    .A(net929),
    .B(net986),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3496_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0358_),
    .B(_0356_),
    .A(_0322_));
 sg13g2_xnor2_1 _3497_ (.Y(_0359_),
    .A(_0321_),
    .B(_0357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3498_ (.Y(_0360_),
    .A(_0355_),
    .B(_0359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3499_ (.B1(_0329_),
    .VDD(VPWR),
    .Y(_0361_),
    .VSS(VGND),
    .A1(_0327_),
    .A2(_0330_));
 sg13g2_nand2_1 _3500_ (.Y(_0362_),
    .A(net931),
    .B(net984),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3501_ (.A(net938),
    .B(net933),
    .C(net981),
    .D(net978),
    .X(_0363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3502_ (.B(net933),
    .C(net981),
    .A(net938),
    .Y(_0364_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net978));
 sg13g2_a22oi_1 _3503_ (.Y(_0365_),
    .B1(net978),
    .B2(net939),
    .A2(net982),
    .A1(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3504_ (.A(_0362_),
    .B(_0363_),
    .C(_0365_),
    .X(_0366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3505_ (.B1(_0362_),
    .VDD(VPWR),
    .Y(_0367_),
    .VSS(VGND),
    .A1(_0363_),
    .A2(_0365_));
 sg13g2_and3_1 _3506_ (.X(_0368_),
    .A(_0361_),
    .B(_0366_),
    .C(_0367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3507_ (.B(_0366_),
    .C(_0367_),
    .A(_0361_),
    .Y(_0369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0366_),
    .A2(_0367_),
    .Y(_0370_),
    .B1(_0361_));
 sg13g2_or3_1 _3509_ (.A(_0360_),
    .B(_0368_),
    .C(_0370_),
    .X(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3510_ (.B1(_0360_),
    .VDD(VPWR),
    .Y(_0372_),
    .VSS(VGND),
    .A1(_0368_),
    .A2(_0370_));
 sg13g2_and3_1 _3511_ (.X(_0373_),
    .A(_0354_),
    .B(_0371_),
    .C(_0372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3512_ (.B(_0371_),
    .C(_0372_),
    .A(_0354_),
    .Y(_0374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3513_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0371_),
    .A2(_0372_),
    .Y(_0375_),
    .B1(_0354_));
 sg13g2_or3_1 _3514_ (.A(_0353_),
    .B(_0373_),
    .C(_0375_),
    .X(_0376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3515_ (.B1(_0353_),
    .VDD(VPWR),
    .Y(_0377_),
    .VSS(VGND),
    .A1(_0373_),
    .A2(_0375_));
 sg13g2_nand3_1 _3516_ (.B(_0376_),
    .C(_0377_),
    .A(_0346_),
    .Y(_0378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3517_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0376_),
    .A2(_0377_),
    .Y(_0379_),
    .B1(_0346_));
 sg13g2_a21o_1 _3518_ (.A2(_0377_),
    .A1(_0376_),
    .B1(_0346_),
    .X(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3519_ (.Y(_0381_),
    .A(_0378_),
    .B(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3520_ (.B(_0381_),
    .A(_0317_),
    .X(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3521_ (.B1(_0343_),
    .VDD(VPWR),
    .Y(_0383_),
    .VSS(VGND),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_nand2_1 _3522_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3523_ (.B(_0383_),
    .A(_0382_),
    .X(_0113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3524_ (.B1(_0374_),
    .VDD(VPWR),
    .Y(_0385_),
    .VSS(VGND),
    .A1(_0353_),
    .A2(_0375_));
 sg13g2_o21ai_1 _3525_ (.B1(_0358_),
    .VDD(VPWR),
    .Y(_0386_),
    .VSS(VGND),
    .A1(_0355_),
    .A2(_0359_));
 sg13g2_nand2_1 _3526_ (.Y(_0387_),
    .A(\DP_1.matrix[0] ),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3527_ (.Y(_0388_),
    .A(net990),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3528_ (.Y(_0389_),
    .A(net990),
    .B(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3529_ (.B(_0389_),
    .A(_0349_),
    .X(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3530_ (.Y(_0391_),
    .B(_0390_),
    .A_N(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3531_ (.Y(_0392_),
    .A(_0387_),
    .B(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3532_ (.Y(_0393_),
    .A(_0386_),
    .B(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3533_ (.Y(_0394_),
    .A(_0386_),
    .B(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3534_ (.Y(_0395_),
    .A(_0350_),
    .B(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3535_ (.B1(_0369_),
    .VDD(VPWR),
    .Y(_0396_),
    .VSS(VGND),
    .A1(_0360_),
    .A2(_0370_));
 sg13g2_nand2_1 _3536_ (.Y(_0397_),
    .A(net988),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3537_ (.Y(_0398_),
    .A(net928),
    .B(net984),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3538_ (.Y(_0399_),
    .A(net929),
    .B(net984),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3539_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0400_),
    .B(_0398_),
    .A(_0357_));
 sg13g2_and2_1 _3540_ (.A(_0356_),
    .B(_0399_),
    .X(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3541_ (.Y(_0402_),
    .A(_0356_),
    .B(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3542_ (.Y(_0403_),
    .A(_0397_),
    .B(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3543_ (.B1(_0364_),
    .VDD(VPWR),
    .Y(_0404_),
    .VSS(VGND),
    .A1(_0362_),
    .A2(_0365_));
 sg13g2_nand2_1 _3544_ (.Y(_0405_),
    .A(net930),
    .B(net981),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3545_ (.A(net938),
    .B(net933),
    .C(net978),
    .D(net1010),
    .X(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3546_ (.B(net934),
    .C(net978),
    .A(net938),
    .Y(_0407_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1010));
 sg13g2_a22oi_1 _3547_ (.Y(_0408_),
    .B1(net1010),
    .B2(net938),
    .A2(net978),
    .A1(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3548_ (.A(_0405_),
    .B(_0406_),
    .C(_0408_),
    .X(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3549_ (.B1(_0405_),
    .VDD(VPWR),
    .Y(_0410_),
    .VSS(VGND),
    .A1(_0406_),
    .A2(_0408_));
 sg13g2_and3_1 _3550_ (.X(_0411_),
    .A(_0404_),
    .B(_0409_),
    .C(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3551_ (.B(_0409_),
    .C(_0410_),
    .A(_0404_),
    .Y(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3552_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0409_),
    .A2(_0410_),
    .Y(_0413_),
    .B1(_0404_));
 sg13g2_or3_1 _3553_ (.A(_0403_),
    .B(_0411_),
    .C(_0413_),
    .X(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3554_ (.B1(_0403_),
    .VDD(VPWR),
    .Y(_0415_),
    .VSS(VGND),
    .A1(_0411_),
    .A2(_0413_));
 sg13g2_and3_1 _3555_ (.X(_0416_),
    .A(_0396_),
    .B(_0414_),
    .C(_0415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3556_ (.B(_0414_),
    .C(_0415_),
    .A(_0396_),
    .Y(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3557_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0414_),
    .A2(_0415_),
    .Y(_0418_),
    .B1(_0396_));
 sg13g2_or3_1 _3558_ (.A(_0395_),
    .B(_0416_),
    .C(_0418_),
    .X(_0419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3559_ (.B1(_0395_),
    .VDD(VPWR),
    .Y(_0420_),
    .VSS(VGND),
    .A1(_0416_),
    .A2(_0418_));
 sg13g2_nand3_1 _3560_ (.B(_0419_),
    .C(_0420_),
    .A(_0385_),
    .Y(_0421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3561_ (.A2(_0420_),
    .A1(_0419_),
    .B1(_0385_),
    .X(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3562_ (.A2(_0422_),
    .A1(_0421_),
    .B1(_0352_),
    .X(_0423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3563_ (.B(_0421_),
    .C(_0422_),
    .A(_0352_),
    .Y(_0424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3564_ (.B1(_0378_),
    .VDD(VPWR),
    .Y(_0425_),
    .VSS(VGND),
    .A1(_0317_),
    .A2(_0379_));
 sg13g2_nand3_1 _3565_ (.B(_0424_),
    .C(_0425_),
    .A(_0423_),
    .Y(_0426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3566_ (.A2(_0424_),
    .A1(_0423_),
    .B1(_0425_),
    .X(_0427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3567_ (.A(_0426_),
    .B(_0427_),
    .X(_0428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3568_ (.B(_0383_),
    .C(_0428_),
    .A(_0382_),
    .Y(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3569_ (.Y(_0114_),
    .A(_0384_),
    .B(_0428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3570_ (.B1(_0393_),
    .VDD(VPWR),
    .Y(_0430_),
    .VSS(VGND),
    .A1(_0350_),
    .A2(_0394_));
 sg13g2_o21ai_1 _3571_ (.B1(_0417_),
    .VDD(VPWR),
    .Y(_0431_),
    .VSS(VGND),
    .A1(_0395_),
    .A2(_0418_));
 sg13g2_o21ai_1 _3572_ (.B1(_0391_),
    .VDD(VPWR),
    .Y(_0432_),
    .VSS(VGND),
    .A1(_0349_),
    .A2(_0389_));
 sg13g2_o21ai_1 _3573_ (.B1(_0400_),
    .VDD(VPWR),
    .Y(_0433_),
    .VSS(VGND),
    .A1(_0397_),
    .A2(_0401_));
 sg13g2_nand2_1 _3574_ (.Y(_0434_),
    .A(net992),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3575_ (.Y(_0435_),
    .A(net988),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3576_ (.Y(_0436_),
    .A(net988),
    .B(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3577_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0437_),
    .B(_0435_),
    .A(_0389_));
 sg13g2_xnor2_1 _3578_ (.Y(_0438_),
    .A(_0388_),
    .B(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3579_ (.B(_0438_),
    .A(_0434_),
    .X(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3580_ (.Y(_0440_),
    .A(_0433_),
    .B(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3581_ (.A(_0440_),
    .B_N(_0432_),
    .Y(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3582_ (.B(_0440_),
    .A(_0432_),
    .X(_0442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3583_ (.B1(_0412_),
    .VDD(VPWR),
    .Y(_0443_),
    .VSS(VGND),
    .A1(_0403_),
    .A2(_0413_));
 sg13g2_nand2_1 _3584_ (.Y(_0444_),
    .A(net986),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3585_ (.Y(_0445_),
    .A(\DP_2.matrix[4] ),
    .B(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3586_ (.Y(_0446_),
    .A(\DP_2.matrix[3] ),
    .B(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3587_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0447_),
    .B(_0445_),
    .A(_0399_));
 sg13g2_and2_1 _3588_ (.A(_0398_),
    .B(_0446_),
    .X(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3589_ (.Y(_0449_),
    .A(_0398_),
    .B(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3590_ (.Y(_0450_),
    .A(_0444_),
    .B(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3591_ (.B1(_0407_),
    .VDD(VPWR),
    .Y(_0451_),
    .VSS(VGND),
    .A1(_0405_),
    .A2(_0408_));
 sg13g2_nand2_1 _3592_ (.Y(_0452_),
    .A(net931),
    .B(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3593_ (.A(net934),
    .B(net930),
    .C(net979),
    .D(net1010),
    .X(_0453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3594_ (.Y(_0454_),
    .B1(net1010),
    .B2(net934),
    .A2(net978),
    .A1(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3595_ (.A(_0453_),
    .B(_0454_),
    .Y(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3596_ (.Y(_0456_),
    .A(_0451_),
    .B(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3597_ (.Y(_0457_),
    .A(_0451_),
    .B(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3598_ (.B(_0457_),
    .A(_0450_),
    .X(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3599_ (.Y(_0459_),
    .A(_0443_),
    .B(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3600_ (.Y(_0460_),
    .A(_0443_),
    .B(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3601_ (.B(_0460_),
    .A(_0442_),
    .X(_0461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3602_ (.Y(_0462_),
    .A(_0431_),
    .B(_0461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3603_ (.Y(_0463_),
    .A(_0431_),
    .B(_0461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3604_ (.Y(_0464_),
    .B(_0430_),
    .A_N(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3605_ (.B(_0463_),
    .A(_0430_),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3606_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0421_),
    .A2(_0424_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_a21o_1 _3607_ (.A2(_0424_),
    .A1(_0421_),
    .B1(_0465_),
    .X(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3608_ (.X(_0468_),
    .A(_0421_),
    .B(_0424_),
    .C(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3609_ (.A(_0466_),
    .B(_0468_),
    .Y(_0469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3610_ (.Y(_0470_),
    .A(_0426_),
    .B(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3611_ (.B(_0470_),
    .A(_0469_),
    .X(_0115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3612_ (.A2(_0439_),
    .A1(_0433_),
    .B1(_0441_),
    .X(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3613_ (.B1(_0459_),
    .VDD(VPWR),
    .Y(_0472_),
    .VSS(VGND),
    .A1(_0442_),
    .A2(_0460_));
 sg13g2_o21ai_1 _3614_ (.B1(_0437_),
    .VDD(VPWR),
    .Y(_0473_),
    .VSS(VGND),
    .A1(_0434_),
    .A2(_0438_));
 sg13g2_o21ai_1 _3615_ (.B1(_0447_),
    .VDD(VPWR),
    .Y(_0474_),
    .VSS(VGND),
    .A1(_0444_),
    .A2(_0448_));
 sg13g2_nand2_1 _3616_ (.Y(_0475_),
    .A(net990),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3617_ (.Y(_0476_),
    .A(net986),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3618_ (.Y(_0477_),
    .A(net986),
    .B(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3619_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0478_),
    .B(_0476_),
    .A(_0436_));
 sg13g2_xnor2_1 _3620_ (.Y(_0479_),
    .A(_0435_),
    .B(_0477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3621_ (.B(_0479_),
    .A(_0475_),
    .X(_0480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3622_ (.Y(_0481_),
    .A(_0474_),
    .B(_0480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3623_ (.A(_0481_),
    .B_N(_0473_),
    .Y(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3624_ (.B(_0481_),
    .A(_0473_),
    .X(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3625_ (.B1(_0456_),
    .VDD(VPWR),
    .Y(_0484_),
    .VSS(VGND),
    .A1(_0450_),
    .A2(_0457_));
 sg13g2_a21oi_1 _3626_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net933),
    .A2(net978),
    .Y(_0485_),
    .B1(_0452_));
 sg13g2_nand2_1 _3627_ (.Y(_0486_),
    .A(net984),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3628_ (.Y(_0487_),
    .A(\DP_2.matrix[4] ),
    .B(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3629_ (.Y(_0488_),
    .A(\DP_2.matrix[3] ),
    .B(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3630_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0489_),
    .B(_0487_),
    .A(_0446_));
 sg13g2_xnor2_1 _3631_ (.Y(_0490_),
    .A(_0445_),
    .B(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3632_ (.B(_0490_),
    .A(_0486_),
    .X(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3633_ (.Y(_0492_),
    .A(_0485_),
    .B(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3634_ (.Y(_0493_),
    .B(_0484_),
    .A_N(_0492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3635_ (.B(_0492_),
    .A(_0484_),
    .X(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3636_ (.B(_0494_),
    .A(_0483_),
    .X(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3637_ (.Y(_0496_),
    .A(_0472_),
    .B(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3638_ (.B(_0495_),
    .A(_0472_),
    .X(_0497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3639_ (.Y(_0498_),
    .A(_0471_),
    .B(_0497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3640_ (.Y(_0499_),
    .A(_0471_),
    .B(_0497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0462_),
    .A2(_0464_),
    .Y(_0500_),
    .B1(_0499_));
 sg13g2_nand3_1 _3642_ (.B(_0464_),
    .C(_0499_),
    .A(_0462_),
    .Y(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3643_ (.A(_0500_),
    .B_N(_0501_),
    .Y(_0502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3644_ (.B(_0383_),
    .C(_0428_),
    .A(_0382_),
    .Y(_0503_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0469_));
 sg13g2_a21oi_1 _3645_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0426_),
    .A2(_0467_),
    .Y(_0504_),
    .B1(_0468_));
 sg13g2_nand2b_1 _3646_ (.Y(_0505_),
    .B(_0503_),
    .A_N(_0504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3647_ (.B(_0505_),
    .A(_0502_),
    .X(_0106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3648_ (.A2(_0480_),
    .A1(_0474_),
    .B1(_0482_),
    .X(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3649_ (.B1(_0493_),
    .VDD(VPWR),
    .Y(_0507_),
    .VSS(VGND),
    .A1(_0483_),
    .A2(_0494_));
 sg13g2_a21o_1 _3650_ (.A2(_0491_),
    .A1(_0485_),
    .B1(_0453_),
    .X(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3651_ (.Y(_0509_),
    .A(\DP_2.matrix[5] ),
    .B(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3652_ (.Y(_0510_),
    .A(\DP_2.matrix[3] ),
    .B(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3653_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0511_),
    .B(_0510_),
    .A(_0487_));
 sg13g2_xnor2_1 _3654_ (.Y(_0512_),
    .A(_0487_),
    .B(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3655_ (.B(_0512_),
    .A(_0509_),
    .X(_0513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3656_ (.Y(_0514_),
    .A(_0508_),
    .B(_0513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3657_ (.B1(_0478_),
    .VDD(VPWR),
    .Y(_0515_),
    .VSS(VGND),
    .A1(_0475_),
    .A2(_0479_));
 sg13g2_inv_1 _3658_ (.VDD(VPWR),
    .Y(_0516_),
    .A(_0515_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3659_ (.B1(_0489_),
    .VDD(VPWR),
    .Y(_0517_),
    .VSS(VGND),
    .A1(_0486_),
    .A2(_0490_));
 sg13g2_nand2_1 _3660_ (.Y(_0518_),
    .A(net988),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3661_ (.Y(_0519_),
    .A(net984),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3662_ (.Y(_0520_),
    .A(net984),
    .B(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3663_ (.B(_0520_),
    .A(_0476_),
    .X(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3664_ (.Y(_0522_),
    .B(_0521_),
    .A_N(_0518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3665_ (.Y(_0523_),
    .A(_0518_),
    .B(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3666_ (.Y(_0524_),
    .A(_0517_),
    .B(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3667_ (.Y(_0525_),
    .A(_0517_),
    .B(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3668_ (.Y(_0526_),
    .A(_0516_),
    .B(_0525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3669_ (.A(_0514_),
    .B(_0526_),
    .Y(_0527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3670_ (.B(_0526_),
    .A(_0514_),
    .X(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3671_ (.Y(_0529_),
    .A(_0507_),
    .B(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3672_ (.A(_0529_),
    .B_N(_0506_),
    .Y(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3673_ (.B(_0529_),
    .A(_0506_),
    .X(_0531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3674_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0496_),
    .A2(_0498_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_nand3_1 _3675_ (.B(_0498_),
    .C(_0531_),
    .A(_0496_),
    .Y(_0533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3676_ (.A(_0532_),
    .B_N(_0533_),
    .Y(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3677_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0502_),
    .A2(_0505_),
    .Y(_0535_),
    .B1(_0500_));
 sg13g2_xnor2_1 _3678_ (.Y(_0107_),
    .A(_0534_),
    .B(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3679_ (.B1(_0524_),
    .VDD(VPWR),
    .Y(_0536_),
    .VSS(VGND),
    .A1(_0516_),
    .A2(_0525_));
 sg13g2_a22oi_1 _3680_ (.Y(_0537_),
    .B1(net1011),
    .B2(\DP_2.matrix[4] ),
    .A2(net980),
    .A1(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3681_ (.Y(_0538_),
    .A(\DP_2.matrix[5] ),
    .B(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3682_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0539_),
    .B(_0538_),
    .A(_0487_));
 sg13g2_nand2b_1 _3683_ (.Y(_0540_),
    .B(_0539_),
    .A_N(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3684_ (.B1(_0522_),
    .VDD(VPWR),
    .Y(_0541_),
    .VSS(VGND),
    .A1(_0476_),
    .A2(_0520_));
 sg13g2_o21ai_1 _3685_ (.B1(_0511_),
    .VDD(VPWR),
    .Y(_0542_),
    .VSS(VGND),
    .A1(_0509_),
    .A2(_0512_));
 sg13g2_nand2_1 _3686_ (.Y(_0543_),
    .A(net986),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3687_ (.Y(_0544_),
    .A(net982),
    .B(\DP_2.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3688_ (.Y(_0545_),
    .A(net982),
    .B(\DP_2.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3689_ (.B(_0545_),
    .A(_0519_),
    .X(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3690_ (.Y(_0547_),
    .B(_0546_),
    .A_N(_0543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3691_ (.Y(_0548_),
    .A(_0543_),
    .B(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3692_ (.Y(_0549_),
    .A(_0542_),
    .B(_0548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3693_ (.A(_0549_),
    .B_N(_0541_),
    .Y(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3694_ (.B(_0549_),
    .A(_0541_),
    .X(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3695_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0552_),
    .B(_0551_),
    .A(_0540_));
 sg13g2_xor2_1 _3696_ (.B(_0551_),
    .A(_0540_),
    .X(_0553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3697_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0508_),
    .A2(_0513_),
    .Y(_0554_),
    .B1(_0527_));
 sg13g2_nor2b_1 _3698_ (.A(_0554_),
    .B_N(_0553_),
    .Y(_0555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3699_ (.Y(_0556_),
    .A(_0553_),
    .B(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3700_ (.Y(_0557_),
    .A(_0536_),
    .B(_0556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0507_),
    .A2(_0528_),
    .Y(_0558_),
    .B1(_0530_));
 sg13g2_nor2_1 _3702_ (.A(_0557_),
    .B(_0558_),
    .Y(_0559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3703_ (.B(_0558_),
    .A(_0557_),
    .X(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3704_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0500_),
    .A2(_0533_),
    .Y(_0561_),
    .B1(_0532_));
 sg13g2_nor2b_1 _3705_ (.A(_0504_),
    .B_N(_0561_),
    .Y(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3706_ (.B1(_0533_),
    .VDD(VPWR),
    .Y(_0563_),
    .VSS(VGND),
    .A1(_0501_),
    .A2(_0532_));
 sg13g2_a21oi_1 _3707_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0503_),
    .A2(_0562_),
    .Y(_0564_),
    .B1(_0563_));
 sg13g2_xor2_1 _3708_ (.B(_0564_),
    .A(_0560_),
    .X(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3709_ (.A2(_0556_),
    .A1(_0536_),
    .B1(_0555_),
    .X(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3710_ (.A2(_0548_),
    .A1(_0542_),
    .B1(_0550_),
    .X(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3711_ (.B1(_0547_),
    .VDD(VPWR),
    .Y(_0567_),
    .VSS(VGND),
    .A1(_0519_),
    .A2(_0545_));
 sg13g2_nand2_1 _3712_ (.Y(_0568_),
    .A(net984),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3713_ (.Y(_0569_),
    .A(net980),
    .B(\DP_2.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3714_ (.Y(_0570_),
    .A(\DP_2.matrix[6] ),
    .B(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3715_ (.B(_0570_),
    .A(_0544_),
    .X(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3716_ (.Y(_0572_),
    .B(_0571_),
    .A_N(_0568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3717_ (.Y(_0573_),
    .A(_0568_),
    .B(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3718_ (.A(_0539_),
    .B_N(_0573_),
    .Y(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3719_ (.Y(_0575_),
    .A(_0539_),
    .B(_0573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3720_ (.Y(_0576_),
    .A(_0567_),
    .B(_0575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3721_ (.A(_0538_),
    .B(_0576_),
    .Y(_0577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3722_ (.B(_0576_),
    .A(_0538_),
    .X(_0578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3723_ (.Y(_0579_),
    .B(_0578_),
    .A_N(_0552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3724_ (.Y(_0580_),
    .A(_0552_),
    .B(_0578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3725_ (.Y(_0581_),
    .A(_0566_),
    .B(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3726_ (.Y(_0582_),
    .A(_0566_),
    .B(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3727_ (.Y(_0583_),
    .B(_0582_),
    .A_N(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3728_ (.A(_0582_),
    .B_N(_0565_),
    .Y(_0584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3729_ (.Y(_0585_),
    .A(_0565_),
    .B(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3730_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0560_),
    .A2(_0564_),
    .Y(_0586_),
    .B1(_0559_));
 sg13g2_xnor2_1 _3731_ (.Y(_0109_),
    .A(_0585_),
    .B(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3732_ (.A(_0560_),
    .B(_0585_),
    .X(_0587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3733_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0564_),
    .C1(_0584_),
    .B1(_0587_),
    .A1(_0559_),
    .Y(_0588_),
    .A2(_0583_));
 sg13g2_and2_1 _3734_ (.A(_0579_),
    .B(_0581_),
    .X(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3735_ (.A2(_0575_),
    .A1(_0567_),
    .B1(_0574_),
    .X(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3736_ (.Y(_0591_),
    .A(net982),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3737_ (.Y(_0592_),
    .A(\DP_2.matrix[7] ),
    .B(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3738_ (.Y(_0593_),
    .A(\DP_2.matrix[6] ),
    .B(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3739_ (.B(_0593_),
    .A(_0569_),
    .X(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3740_ (.Y(_0595_),
    .B(_0594_),
    .A_N(_0591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3741_ (.Y(_0596_),
    .A(_0591_),
    .B(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3742_ (.B1(_0572_),
    .VDD(VPWR),
    .Y(_0597_),
    .VSS(VGND),
    .A1(_0544_),
    .A2(_0570_));
 sg13g2_nand2_1 _3743_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3744_ (.B(_0597_),
    .A(_0596_),
    .X(_0599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3745_ (.Y(_0600_),
    .A(_0577_),
    .B(_0599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3746_ (.A(_0600_),
    .B_N(_0590_),
    .Y(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3747_ (.B(_0600_),
    .A(_0590_),
    .X(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3748_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0603_),
    .B(_0602_),
    .A(_0589_));
 sg13g2_xor2_1 _3749_ (.B(_0602_),
    .A(_0589_),
    .X(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3750_ (.VDD(VPWR),
    .Y(_0605_),
    .A(_0604_),
    .VSS(VGND));
 sg13g2_xnor2_1 _3751_ (.Y(_0110_),
    .A(_0588_),
    .B(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3752_ (.B1(_0603_),
    .VDD(VPWR),
    .Y(_0606_),
    .VSS(VGND),
    .A1(_0588_),
    .A2(_0605_));
 sg13g2_a21oi_1 _3753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0577_),
    .A2(_0599_),
    .Y(_0607_),
    .B1(_0601_));
 sg13g2_o21ai_1 _3754_ (.B1(_0595_),
    .VDD(VPWR),
    .Y(_0608_),
    .VSS(VGND),
    .A1(_0569_),
    .A2(_0593_));
 sg13g2_nand2_1 _3755_ (.Y(_0609_),
    .A(net980),
    .B(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3756_ (.B(_0609_),
    .A(_0592_),
    .X(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3757_ (.Y(_0611_),
    .A(_0608_),
    .B(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3758_ (.Y(_0612_),
    .A(_0598_),
    .B(_0611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3759_ (.Y(_0613_),
    .A(_0607_),
    .B(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3760_ (.Y(_0111_),
    .A(_0606_),
    .B(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3761_ (.A(net977),
    .B(net924),
    .X(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3762_ (.X(_0614_),
    .A(net975),
    .B(net918),
    .C(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3763_ (.Y(_0615_),
    .B1(net918),
    .B2(net977),
    .A2(net975),
    .A1(net924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3764_ (.A(_0614_),
    .B(_0615_),
    .Y(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3765_ (.A(net977),
    .B(net916),
    .X(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3766_ (.A(net924),
    .B(net975),
    .C(net918),
    .D(net973),
    .X(_0617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3767_ (.Y(_0618_),
    .B1(net973),
    .B2(net924),
    .A2(net918),
    .A1(net975),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3768_ (.A(_0617_),
    .B(_0618_),
    .Y(_0619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3769_ (.B(_0619_),
    .A(_0616_),
    .X(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3770_ (.Y(_0621_),
    .A(_0614_),
    .B(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3771_ (.B(_0620_),
    .A(_0614_),
    .X(_0076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3772_ (.Y(_0622_),
    .A(net281),
    .B(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0616_),
    .A2(_0619_),
    .Y(_0623_),
    .B1(_0617_));
 sg13g2_nand2_1 _3774_ (.Y(_0624_),
    .A(net975),
    .B(net916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3775_ (.A(net924),
    .B(net918),
    .C(net973),
    .D(net972),
    .X(_0625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3776_ (.B(net918),
    .C(net973),
    .A(net924),
    .Y(_0626_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net972));
 sg13g2_a22oi_1 _3777_ (.Y(_0627_),
    .B1(net972),
    .B2(net924),
    .A2(net973),
    .A1(net918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3778_ (.A(_0624_),
    .B(_0625_),
    .C(_0627_),
    .Y(_0628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3779_ (.B1(_0624_),
    .VDD(VPWR),
    .Y(_0629_),
    .VSS(VGND),
    .A1(_0625_),
    .A2(_0627_));
 sg13g2_nor2b_1 _3780_ (.A(_0628_),
    .B_N(_0629_),
    .Y(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3781_ (.Y(_0631_),
    .B(_0630_),
    .A_N(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3782_ (.Y(_0632_),
    .A(_0623_),
    .B(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3783_ (.Y(_0633_),
    .B(_0632_),
    .A_N(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3784_ (.Y(_0634_),
    .A(_0622_),
    .B(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3785_ (.A(_0621_),
    .B_N(_0634_),
    .Y(_0635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3786_ (.Y(_0077_),
    .A(_0621_),
    .B(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3787_ (.Y(_0636_),
    .B1(\DP_2.matrix[40] ),
    .B2(net977),
    .A2(net915),
    .A1(net975),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3788_ (.Y(_0637_),
    .A(net975),
    .B(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3789_ (.A(_0622_),
    .B(_0637_),
    .Y(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3790_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0639_),
    .B(_0638_),
    .A(_0636_));
 sg13g2_o21ai_1 _3791_ (.B1(_0626_),
    .VDD(VPWR),
    .Y(_0640_),
    .VSS(VGND),
    .A1(_0624_),
    .A2(_0627_));
 sg13g2_nand2_1 _3792_ (.Y(_0641_),
    .A(net973),
    .B(net916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3793_ (.A(net923),
    .B(\DP_2.matrix[37] ),
    .C(net972),
    .D(net970),
    .X(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3794_ (.B(net921),
    .C(net971),
    .A(net923),
    .Y(_0643_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net970));
 sg13g2_a22oi_1 _3795_ (.Y(_0644_),
    .B1(net970),
    .B2(net923),
    .A2(net971),
    .A1(net921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3796_ (.A(_0641_),
    .B(_0642_),
    .C(_0644_),
    .X(_0645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3797_ (.B1(_0641_),
    .VDD(VPWR),
    .Y(_0646_),
    .VSS(VGND),
    .A1(_0642_),
    .A2(_0644_));
 sg13g2_nand3_1 _3798_ (.B(_0645_),
    .C(_0646_),
    .A(_0640_),
    .Y(_0647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3799_ (.A2(_0646_),
    .A1(_0645_),
    .B1(_0640_),
    .X(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3800_ (.Y(_0649_),
    .A(_0647_),
    .B(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3801_ (.B(_0649_),
    .A(_0639_),
    .X(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3802_ (.Y(_0651_),
    .A(_0631_),
    .B(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3803_ (.Y(_0652_),
    .A(_0650_),
    .B(_0651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3804_ (.B(_0651_),
    .A(_0650_),
    .X(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3805_ (.A(_0635_),
    .B(_0653_),
    .X(_0654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3806_ (.B(_0653_),
    .A(_0635_),
    .X(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3807_ (.B1(_0647_),
    .VDD(VPWR),
    .Y(_0655_),
    .VSS(VGND),
    .A1(_0639_),
    .A2(_0649_));
 sg13g2_nand2_1 _3808_ (.Y(_0656_),
    .A(net977),
    .B(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3809_ (.Y(_0657_),
    .A(net974),
    .B(net912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3810_ (.Y(_0658_),
    .A(net974),
    .B(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3811_ (.B(_0658_),
    .A(_0637_),
    .X(_0659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3812_ (.Y(_0660_),
    .B(_0659_),
    .A_N(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3813_ (.B(_0659_),
    .A(_0656_),
    .X(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3814_ (.B1(_0643_),
    .VDD(VPWR),
    .Y(_0662_),
    .VSS(VGND),
    .A1(_0641_),
    .A2(_0644_));
 sg13g2_nand2_1 _3815_ (.Y(_0663_),
    .A(net917),
    .B(net971),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3816_ (.A(net923),
    .B(net921),
    .C(net969),
    .D(\DP_1.matrix[41] ),
    .X(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3817_ (.B(net921),
    .C(net969),
    .A(net923),
    .Y(_0665_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net967));
 sg13g2_a22oi_1 _3818_ (.Y(_0666_),
    .B1(net967),
    .B2(net923),
    .A2(net969),
    .A1(net921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3819_ (.A(_0663_),
    .B(_0664_),
    .C(_0666_),
    .X(_0667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3820_ (.B1(_0663_),
    .VDD(VPWR),
    .Y(_0668_),
    .VSS(VGND),
    .A1(_0664_),
    .A2(_0666_));
 sg13g2_and3_1 _3821_ (.X(_0669_),
    .A(_0662_),
    .B(_0667_),
    .C(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3822_ (.B(_0667_),
    .C(_0668_),
    .A(_0662_),
    .Y(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0667_),
    .A2(_0668_),
    .Y(_0671_),
    .B1(_0662_));
 sg13g2_or3_1 _3824_ (.A(_0661_),
    .B(_0669_),
    .C(_0671_),
    .X(_0672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3825_ (.B1(_0661_),
    .VDD(VPWR),
    .Y(_0673_),
    .VSS(VGND),
    .A1(_0669_),
    .A2(_0671_));
 sg13g2_nand3_1 _3826_ (.B(_0672_),
    .C(_0673_),
    .A(_0655_),
    .Y(_0674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3827_ (.A2(_0673_),
    .A1(_0672_),
    .B1(_0655_),
    .X(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3828_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0674_),
    .A2(_0675_),
    .Y(_0676_),
    .B1(_0638_));
 sg13g2_and3_1 _3829_ (.X(_0677_),
    .A(_0638_),
    .B(_0674_),
    .C(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3830_ (.B(_0674_),
    .C(_0675_),
    .A(_0638_),
    .Y(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3831_ (.A(_0652_),
    .B(_0676_),
    .C(_0677_),
    .Y(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3832_ (.B1(_0652_),
    .VDD(VPWR),
    .Y(_0680_),
    .VSS(VGND),
    .A1(_0676_),
    .A2(_0677_));
 sg13g2_nand2b_1 _3833_ (.Y(_0681_),
    .B(_0680_),
    .A_N(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3834_ (.Y(_0116_),
    .A(_0654_),
    .B(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3835_ (.Y(_0682_),
    .A(_0674_),
    .B(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3836_ (.B1(_0660_),
    .VDD(VPWR),
    .Y(_0683_),
    .VSS(VGND),
    .A1(_0637_),
    .A2(_0658_));
 sg13g2_nand2_1 _3837_ (.Y(_0684_),
    .A(net977),
    .B(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3838_ (.Y(_0685_),
    .B(_0683_),
    .A_N(_0684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3839_ (.B(_0684_),
    .A(_0683_),
    .X(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3840_ (.B1(_0670_),
    .VDD(VPWR),
    .Y(_0687_),
    .VSS(VGND),
    .A1(_0661_),
    .A2(_0671_));
 sg13g2_nand2_1 _3841_ (.Y(_0688_),
    .A(net976),
    .B(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3842_ (.Y(_0689_),
    .A(net972),
    .B(net912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3843_ (.Y(_0690_),
    .A(net972),
    .B(net914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3844_ (.B(_0690_),
    .A(_0657_),
    .X(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3845_ (.Y(_0692_),
    .B(_0691_),
    .A_N(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3846_ (.Y(_0693_),
    .A(_0688_),
    .B(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3847_ (.B1(_0665_),
    .VDD(VPWR),
    .Y(_0694_),
    .VSS(VGND),
    .A1(_0663_),
    .A2(_0666_));
 sg13g2_nand2_1 _3848_ (.Y(_0695_),
    .A(net917),
    .B(net968),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3849_ (.A(net922),
    .B(net921),
    .C(net967),
    .D(net965),
    .X(_0696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3850_ (.B(net920),
    .C(net967),
    .A(net922),
    .Y(_0697_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net965));
 sg13g2_a22oi_1 _3851_ (.Y(_0698_),
    .B1(net965),
    .B2(net922),
    .A2(net967),
    .A1(net920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3852_ (.A(_0695_),
    .B(_0696_),
    .C(_0698_),
    .X(_0699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3853_ (.B1(_0695_),
    .VDD(VPWR),
    .Y(_0700_),
    .VSS(VGND),
    .A1(_0696_),
    .A2(_0698_));
 sg13g2_and3_1 _3854_ (.X(_0701_),
    .A(_0694_),
    .B(_0699_),
    .C(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3855_ (.B(_0699_),
    .C(_0700_),
    .A(_0694_),
    .Y(_0702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3856_ (.A2(_0700_),
    .A1(_0699_),
    .B1(_0694_),
    .X(_0703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3857_ (.B(_0702_),
    .C(_0703_),
    .A(_0693_),
    .Y(_0704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3858_ (.A2(_0703_),
    .A1(_0702_),
    .B1(_0693_),
    .X(_0705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3859_ (.B(_0704_),
    .C(_0705_),
    .A(_0687_),
    .Y(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0704_),
    .A2(_0705_),
    .Y(_0707_),
    .B1(_0687_));
 sg13g2_a21o_1 _3861_ (.A2(_0705_),
    .A1(_0704_),
    .B1(_0687_),
    .X(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3862_ (.Y(_0709_),
    .A(_0706_),
    .B(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3863_ (.Y(_0710_),
    .A(_0686_),
    .B(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3864_ (.Y(_0711_),
    .B(_0682_),
    .A_N(_0710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3865_ (.B(_0710_),
    .A(_0682_),
    .X(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0654_),
    .A2(_0680_),
    .Y(_0713_),
    .B1(_0679_));
 sg13g2_xor2_1 _3867_ (.B(_0713_),
    .A(_0712_),
    .X(_0123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3868_ (.B1(_0706_),
    .VDD(VPWR),
    .Y(_0714_),
    .VSS(VGND),
    .A1(_0686_),
    .A2(_0707_));
 sg13g2_o21ai_1 _3869_ (.B1(_0692_),
    .VDD(VPWR),
    .Y(_0715_),
    .VSS(VGND),
    .A1(_0657_),
    .A2(_0690_));
 sg13g2_a22oi_1 _3870_ (.Y(_0716_),
    .B1(net906),
    .B2(\DP_1.matrix[36] ),
    .A2(net908),
    .A1(net976),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3871_ (.Y(_0717_),
    .A(net976),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3872_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0718_),
    .B(_0717_),
    .A(_0684_));
 sg13g2_nor2b_1 _3873_ (.A(_0716_),
    .B_N(_0718_),
    .Y(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3874_ (.A(_0715_),
    .B(_0719_),
    .X(_0720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3875_ (.Y(_0721_),
    .A(_0715_),
    .B(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3876_ (.A2(_0703_),
    .A1(_0693_),
    .B1(_0701_),
    .X(_0722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3877_ (.Y(_0723_),
    .A(net973),
    .B(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3878_ (.Y(_0724_),
    .A(net914),
    .B(net968),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3879_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0725_),
    .B(_0724_),
    .A(_0689_));
 sg13g2_xnor2_1 _3880_ (.Y(_0726_),
    .A(_0689_),
    .B(_0724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3881_ (.Y(_0727_),
    .A(_0723_),
    .B(_0726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3882_ (.B1(_0697_),
    .VDD(VPWR),
    .Y(_0728_),
    .VSS(VGND),
    .A1(_0695_),
    .A2(_0698_));
 sg13g2_nand2_1 _3883_ (.Y(_0729_),
    .A(net916),
    .B(net966),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3884_ (.A(\DP_2.matrix[36] ),
    .B(net919),
    .C(net963),
    .D(net962),
    .X(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3885_ (.B(net919),
    .C(net963),
    .A(net922),
    .Y(_0731_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net960));
 sg13g2_a22oi_1 _3886_ (.Y(_0732_),
    .B1(net960),
    .B2(net922),
    .A2(net963),
    .A1(net919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3887_ (.A(_0729_),
    .B(_0730_),
    .C(_0732_),
    .X(_0733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3888_ (.B1(_0729_),
    .VDD(VPWR),
    .Y(_0734_),
    .VSS(VGND),
    .A1(_0730_),
    .A2(_0732_));
 sg13g2_and3_1 _3889_ (.X(_0735_),
    .A(_0728_),
    .B(_0733_),
    .C(_0734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3890_ (.B(_0733_),
    .C(_0734_),
    .A(_0728_),
    .Y(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3891_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0733_),
    .A2(_0734_),
    .Y(_0737_),
    .B1(_0728_));
 sg13g2_or3_1 _3892_ (.A(_0727_),
    .B(_0735_),
    .C(_0737_),
    .X(_0738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3893_ (.B1(_0727_),
    .VDD(VPWR),
    .Y(_0739_),
    .VSS(VGND),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_and3_1 _3894_ (.X(_0740_),
    .A(_0722_),
    .B(_0738_),
    .C(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3895_ (.B(_0738_),
    .C(_0739_),
    .A(_0722_),
    .Y(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3896_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0738_),
    .A2(_0739_),
    .Y(_0742_),
    .B1(_0722_));
 sg13g2_or3_1 _3897_ (.A(_0721_),
    .B(_0740_),
    .C(_0742_),
    .X(_0743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3898_ (.B1(_0721_),
    .VDD(VPWR),
    .Y(_0744_),
    .VSS(VGND),
    .A1(_0740_),
    .A2(_0742_));
 sg13g2_nand3_1 _3899_ (.B(_0743_),
    .C(_0744_),
    .A(_0714_),
    .Y(_0745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3900_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0743_),
    .A2(_0744_),
    .Y(_0746_),
    .B1(_0714_));
 sg13g2_a21o_1 _3901_ (.A2(_0744_),
    .A1(_0743_),
    .B1(_0714_),
    .X(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3902_ (.Y(_0748_),
    .A(_0745_),
    .B(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3903_ (.B(_0748_),
    .A(_0685_),
    .X(_0749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3904_ (.B1(_0711_),
    .VDD(VPWR),
    .Y(_0750_),
    .VSS(VGND),
    .A1(_0712_),
    .A2(_0713_));
 sg13g2_nand2_1 _3905_ (.Y(_0751_),
    .A(_0749_),
    .B(_0750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3906_ (.B(_0750_),
    .A(_0749_),
    .X(_0124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3907_ (.B1(_0741_),
    .VDD(VPWR),
    .Y(_0752_),
    .VSS(VGND),
    .A1(_0721_),
    .A2(_0742_));
 sg13g2_o21ai_1 _3908_ (.B1(_0725_),
    .VDD(VPWR),
    .Y(_0753_),
    .VSS(VGND),
    .A1(_0723_),
    .A2(_0726_));
 sg13g2_nand2_1 _3909_ (.Y(_0754_),
    .A(net977),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3910_ (.Y(_0755_),
    .A(net974),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3911_ (.Y(_0756_),
    .A(net974),
    .B(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3912_ (.B(_0756_),
    .A(_0717_),
    .X(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3913_ (.Y(_0758_),
    .B(_0757_),
    .A_N(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3914_ (.Y(_0759_),
    .A(_0754_),
    .B(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3915_ (.Y(_0760_),
    .A(_0753_),
    .B(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3916_ (.Y(_0761_),
    .A(_0753_),
    .B(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3917_ (.Y(_0762_),
    .A(_0718_),
    .B(_0761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3918_ (.B1(_0736_),
    .VDD(VPWR),
    .Y(_0763_),
    .VSS(VGND),
    .A1(_0727_),
    .A2(_0737_));
 sg13g2_nand2_1 _3919_ (.Y(_0764_),
    .A(net971),
    .B(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3920_ (.Y(_0765_),
    .A(net912),
    .B(net967),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3921_ (.A(net914),
    .B(net968),
    .C(net912),
    .D(net966),
    .X(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3922_ (.Y(_0767_),
    .B1(net966),
    .B2(net914),
    .A2(net912),
    .A1(net969),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3923_ (.A(_0764_),
    .B(_0766_),
    .C(_0767_),
    .Y(_0768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3924_ (.B1(_0764_),
    .VDD(VPWR),
    .Y(_0769_),
    .VSS(VGND),
    .A1(_0766_),
    .A2(_0767_));
 sg13g2_nand2b_1 _3925_ (.Y(_0770_),
    .B(_0769_),
    .A_N(_0768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3926_ (.B1(_0731_),
    .VDD(VPWR),
    .Y(_0771_),
    .VSS(VGND),
    .A1(_0729_),
    .A2(_0732_));
 sg13g2_nand2_1 _3927_ (.Y(_0772_),
    .A(net916),
    .B(net963),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3928_ (.A(net922),
    .B(net919),
    .C(net960),
    .D(net1008),
    .X(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3929_ (.B(net919),
    .C(net960),
    .A(net922),
    .Y(_0774_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1008));
 sg13g2_a22oi_1 _3930_ (.Y(_0775_),
    .B1(net1008),
    .B2(net922),
    .A2(net960),
    .A1(net920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3931_ (.A(_0772_),
    .B(_0773_),
    .C(_0775_),
    .X(_0776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3932_ (.B1(_0772_),
    .VDD(VPWR),
    .Y(_0777_),
    .VSS(VGND),
    .A1(_0773_),
    .A2(_0775_));
 sg13g2_and3_1 _3933_ (.X(_0778_),
    .A(_0771_),
    .B(_0776_),
    .C(_0777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3934_ (.B(_0776_),
    .C(_0777_),
    .A(_0771_),
    .Y(_0779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3935_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0776_),
    .A2(_0777_),
    .Y(_0780_),
    .B1(_0771_));
 sg13g2_or3_1 _3936_ (.A(_0770_),
    .B(_0778_),
    .C(_0780_),
    .X(_0781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3937_ (.B1(_0770_),
    .VDD(VPWR),
    .Y(_0782_),
    .VSS(VGND),
    .A1(_0778_),
    .A2(_0780_));
 sg13g2_and3_1 _3938_ (.X(_0783_),
    .A(_0763_),
    .B(_0781_),
    .C(_0782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3939_ (.B(_0781_),
    .C(_0782_),
    .A(_0763_),
    .Y(_0784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0781_),
    .A2(_0782_),
    .Y(_0785_),
    .B1(_0763_));
 sg13g2_or3_1 _3941_ (.A(_0762_),
    .B(_0783_),
    .C(_0785_),
    .X(_0786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3942_ (.B1(_0762_),
    .VDD(VPWR),
    .Y(_0787_),
    .VSS(VGND),
    .A1(_0783_),
    .A2(_0785_));
 sg13g2_nand3_1 _3943_ (.B(_0786_),
    .C(_0787_),
    .A(_0752_),
    .Y(_0788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3944_ (.A2(_0787_),
    .A1(_0786_),
    .B1(_0752_),
    .X(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3945_ (.A2(_0789_),
    .A1(_0788_),
    .B1(_0720_),
    .X(_0790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3946_ (.B(_0788_),
    .C(_0789_),
    .A(_0720_),
    .Y(_0791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3947_ (.B1(_0745_),
    .VDD(VPWR),
    .Y(_0792_),
    .VSS(VGND),
    .A1(_0685_),
    .A2(_0746_));
 sg13g2_nand3_1 _3948_ (.B(_0791_),
    .C(_0792_),
    .A(_0790_),
    .Y(_0793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3949_ (.A2(_0791_),
    .A1(_0790_),
    .B1(_0792_),
    .X(_0794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3950_ (.A(_0793_),
    .B(_0794_),
    .X(_0795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3951_ (.B(_0750_),
    .C(_0795_),
    .A(_0749_),
    .Y(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3952_ (.Y(_0125_),
    .A(_0751_),
    .B(_0795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3953_ (.B1(_0760_),
    .VDD(VPWR),
    .Y(_0797_),
    .VSS(VGND),
    .A1(_0718_),
    .A2(_0761_));
 sg13g2_o21ai_1 _3954_ (.B1(_0784_),
    .VDD(VPWR),
    .Y(_0798_),
    .VSS(VGND),
    .A1(_0762_),
    .A2(_0785_));
 sg13g2_o21ai_1 _3955_ (.B1(_0758_),
    .VDD(VPWR),
    .Y(_0799_),
    .VSS(VGND),
    .A1(_0717_),
    .A2(_0756_));
 sg13g2_or2_1 _3956_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0800_),
    .B(_0768_),
    .A(_0766_));
 sg13g2_nand2_1 _3957_ (.Y(_0801_),
    .A(net976),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3958_ (.Y(_0802_),
    .A(net971),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3959_ (.Y(_0803_),
    .A(net971),
    .B(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3960_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0804_),
    .B(_0802_),
    .A(_0756_));
 sg13g2_xnor2_1 _3961_ (.Y(_0805_),
    .A(_0755_),
    .B(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3962_ (.B(_0805_),
    .A(_0801_),
    .X(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3963_ (.Y(_0807_),
    .A(_0800_),
    .B(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3964_ (.A(_0807_),
    .B_N(_0799_),
    .Y(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3965_ (.B(_0807_),
    .A(_0799_),
    .X(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3966_ (.B1(_0779_),
    .VDD(VPWR),
    .Y(_0810_),
    .VSS(VGND),
    .A1(_0770_),
    .A2(_0780_));
 sg13g2_nand2_1 _3967_ (.Y(_0811_),
    .A(net968),
    .B(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3968_ (.Y(_0812_),
    .A(net914),
    .B(net963),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3969_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0813_),
    .B(_0812_),
    .A(_0765_));
 sg13g2_and2_1 _3970_ (.A(_0765_),
    .B(_0812_),
    .X(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3971_ (.Y(_0815_),
    .A(_0765_),
    .B(_0812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3972_ (.Y(_0816_),
    .A(_0811_),
    .B(_0815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3973_ (.B1(_0774_),
    .VDD(VPWR),
    .Y(_0817_),
    .VSS(VGND),
    .A1(_0772_),
    .A2(_0775_));
 sg13g2_nand2_1 _3974_ (.Y(_0818_),
    .A(net916),
    .B(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3975_ (.A(net919),
    .B(net917),
    .C(net960),
    .D(net1008),
    .X(_0819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3976_ (.Y(_0820_),
    .B1(net1008),
    .B2(net919),
    .A2(net960),
    .A1(net917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3977_ (.A(_0819_),
    .B(_0820_),
    .Y(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3978_ (.Y(_0822_),
    .A(_0817_),
    .B(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3979_ (.Y(_0823_),
    .A(_0817_),
    .B(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3980_ (.B(_0823_),
    .A(_0816_),
    .X(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3981_ (.Y(_0825_),
    .A(_0810_),
    .B(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3982_ (.Y(_0826_),
    .A(_0810_),
    .B(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3983_ (.B(_0826_),
    .A(_0809_),
    .X(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3984_ (.Y(_0828_),
    .A(_0798_),
    .B(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3985_ (.Y(_0829_),
    .A(_0798_),
    .B(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3986_ (.Y(_0830_),
    .B(_0797_),
    .A_N(_0829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3987_ (.B(_0829_),
    .A(_0797_),
    .X(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3988_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0788_),
    .A2(_0791_),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_a21o_1 _3989_ (.A2(_0791_),
    .A1(_0788_),
    .B1(_0831_),
    .X(_0833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3990_ (.X(_0834_),
    .A(_0788_),
    .B(_0791_),
    .C(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3991_ (.A(_0832_),
    .B(_0834_),
    .Y(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3992_ (.Y(_0836_),
    .A(_0793_),
    .B(_0796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3993_ (.B(_0836_),
    .A(_0835_),
    .X(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3994_ (.A2(_0806_),
    .A1(_0800_),
    .B1(_0808_),
    .X(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3995_ (.B1(_0825_),
    .VDD(VPWR),
    .Y(_0838_),
    .VSS(VGND),
    .A1(_0809_),
    .A2(_0826_));
 sg13g2_o21ai_1 _3996_ (.B1(_0804_),
    .VDD(VPWR),
    .Y(_0839_),
    .VSS(VGND),
    .A1(_0801_),
    .A2(_0805_));
 sg13g2_o21ai_1 _3997_ (.B1(_0813_),
    .VDD(VPWR),
    .Y(_0840_),
    .VSS(VGND),
    .A1(_0811_),
    .A2(_0814_));
 sg13g2_nand2_1 _3998_ (.Y(_0841_),
    .A(net974),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3999_ (.Y(_0842_),
    .A(net968),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4000_ (.Y(_0843_),
    .A(net968),
    .B(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4001_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0844_),
    .B(_0842_),
    .A(_0803_));
 sg13g2_xnor2_1 _4002_ (.Y(_0845_),
    .A(_0802_),
    .B(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4003_ (.B(_0845_),
    .A(_0841_),
    .X(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4004_ (.Y(_0847_),
    .A(_0840_),
    .B(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4005_ (.A(_0847_),
    .B_N(_0839_),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4006_ (.B(_0847_),
    .A(_0839_),
    .X(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4007_ (.B1(_0822_),
    .VDD(VPWR),
    .Y(_0850_),
    .VSS(VGND),
    .A1(_0816_),
    .A2(_0823_));
 sg13g2_a21oi_1 _4008_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net919),
    .A2(net960),
    .Y(_0851_),
    .B1(_0818_));
 sg13g2_nand2_1 _4009_ (.Y(_0852_),
    .A(net966),
    .B(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4010_ (.Y(_0853_),
    .A(net912),
    .B(net961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4011_ (.A(net914),
    .B(net912),
    .C(net963),
    .D(net961),
    .X(_0854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4012_ (.Y(_0855_),
    .B1(net961),
    .B2(net914),
    .A2(net963),
    .A1(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4013_ (.A(_0852_),
    .B(_0854_),
    .C(_0855_),
    .Y(_0856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4014_ (.B1(_0852_),
    .VDD(VPWR),
    .Y(_0857_),
    .VSS(VGND),
    .A1(_0854_),
    .A2(_0855_));
 sg13g2_nor2b_1 _4015_ (.A(_0856_),
    .B_N(_0857_),
    .Y(_0858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4016_ (.Y(_0859_),
    .A(_0851_),
    .B(_0858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4017_ (.Y(_0860_),
    .B(_0850_),
    .A_N(_0859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4018_ (.B(_0859_),
    .A(_0850_),
    .X(_0861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4019_ (.B(_0861_),
    .A(_0849_),
    .X(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4020_ (.Y(_0863_),
    .A(_0838_),
    .B(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4021_ (.B(_0862_),
    .A(_0838_),
    .X(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4022_ (.Y(_0865_),
    .A(_0837_),
    .B(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4023_ (.Y(_0866_),
    .A(_0837_),
    .B(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4024_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0828_),
    .A2(_0830_),
    .Y(_0867_),
    .B1(_0866_));
 sg13g2_nand3_1 _4025_ (.B(_0830_),
    .C(_0866_),
    .A(_0828_),
    .Y(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4026_ (.A(_0867_),
    .B_N(_0868_),
    .Y(_0869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4027_ (.B(_0750_),
    .C(_0795_),
    .A(_0749_),
    .Y(_0870_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0835_));
 sg13g2_a21oi_1 _4028_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0793_),
    .A2(_0833_),
    .Y(_0871_),
    .B1(_0834_));
 sg13g2_nand2b_1 _4029_ (.Y(_0872_),
    .B(_0870_),
    .A_N(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4030_ (.B(_0872_),
    .A(_0869_),
    .X(_0117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4031_ (.A2(_0846_),
    .A1(_0840_),
    .B1(_0848_),
    .X(_0873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4032_ (.B1(_0860_),
    .VDD(VPWR),
    .Y(_0874_),
    .VSS(VGND),
    .A1(_0849_),
    .A2(_0861_));
 sg13g2_a21o_1 _4033_ (.A2(_0858_),
    .A1(_0851_),
    .B1(_0819_),
    .X(_0875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4034_ (.Y(_0876_),
    .A(net910),
    .B(net964),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4035_ (.Y(_0877_),
    .A(net915),
    .B(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4036_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0878_),
    .B(_0877_),
    .A(_0853_));
 sg13g2_xnor2_1 _4037_ (.Y(_0879_),
    .A(_0853_),
    .B(_0877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4038_ (.B(_0879_),
    .A(_0876_),
    .X(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4039_ (.Y(_0881_),
    .A(_0875_),
    .B(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4040_ (.B1(_0844_),
    .VDD(VPWR),
    .Y(_0882_),
    .VSS(VGND),
    .A1(_0841_),
    .A2(_0845_));
 sg13g2_or2_1 _4041_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0883_),
    .B(_0856_),
    .A(_0854_));
 sg13g2_nand2_1 _4042_ (.Y(_0884_),
    .A(net971),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4043_ (.Y(_0885_),
    .A(net966),
    .B(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4044_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0886_),
    .B(_0885_),
    .A(_0842_));
 sg13g2_xnor2_1 _4045_ (.Y(_0887_),
    .A(_0842_),
    .B(_0885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4046_ (.B(_0887_),
    .A(_0884_),
    .X(_0888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4047_ (.Y(_0889_),
    .A(_0883_),
    .B(_0888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4048_ (.A(_0889_),
    .B_N(_0882_),
    .Y(_0890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4049_ (.B(_0889_),
    .A(_0882_),
    .X(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4050_ (.A(_0881_),
    .B(_0891_),
    .Y(_0892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4051_ (.B(_0891_),
    .A(_0881_),
    .X(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4052_ (.Y(_0894_),
    .A(_0874_),
    .B(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4053_ (.A(_0894_),
    .B_N(_0873_),
    .Y(_0895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4054_ (.B(_0894_),
    .A(_0873_),
    .X(_0896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4055_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0863_),
    .A2(_0865_),
    .Y(_0897_),
    .B1(_0896_));
 sg13g2_nand3_1 _4056_ (.B(_0865_),
    .C(_0896_),
    .A(_0863_),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4057_ (.A(_0897_),
    .B_N(_0898_),
    .Y(_0899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4058_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0869_),
    .A2(_0872_),
    .Y(_0900_),
    .B1(_0867_));
 sg13g2_xnor2_1 _4059_ (.Y(_0118_),
    .A(_0899_),
    .B(_0900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4060_ (.A2(_0888_),
    .A1(_0883_),
    .B1(_0890_),
    .X(_0901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4061_ (.Y(_0902_),
    .B1(net1009),
    .B2(net913),
    .A2(net961),
    .A1(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4062_ (.Y(_0903_),
    .A(net910),
    .B(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4063_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0904_),
    .B(_0903_),
    .A(_0853_));
 sg13g2_nand2b_1 _4064_ (.Y(_0905_),
    .B(_0904_),
    .A_N(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4065_ (.B1(_0886_),
    .VDD(VPWR),
    .Y(_0906_),
    .VSS(VGND),
    .A1(_0884_),
    .A2(_0887_));
 sg13g2_o21ai_1 _4066_ (.B1(_0878_),
    .VDD(VPWR),
    .Y(_0907_),
    .VSS(VGND),
    .A1(_0876_),
    .A2(_0879_));
 sg13g2_nand2_1 _4067_ (.Y(_0908_),
    .A(net968),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4068_ (.Y(_0909_),
    .A(net964),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4069_ (.A(_0885_),
    .B(_0909_),
    .Y(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4070_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0911_),
    .B(_0909_),
    .A(_0885_));
 sg13g2_a22oi_1 _4071_ (.Y(_0912_),
    .B1(net906),
    .B2(net966),
    .A2(net908),
    .A1(net964),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4072_ (.A(_0910_),
    .B(_0912_),
    .Y(_0913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4073_ (.Y(_0914_),
    .A(_0908_),
    .B(_0913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4074_ (.Y(_0915_),
    .A(_0907_),
    .B(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4075_ (.A(_0915_),
    .B_N(_0906_),
    .Y(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4076_ (.B(_0915_),
    .A(_0906_),
    .X(_0917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4077_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0918_),
    .B(_0917_),
    .A(_0905_));
 sg13g2_xor2_1 _4078_ (.B(_0917_),
    .A(_0905_),
    .X(_0919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4079_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0875_),
    .A2(_0880_),
    .Y(_0920_),
    .B1(_0892_));
 sg13g2_nor2b_1 _4080_ (.A(_0920_),
    .B_N(_0919_),
    .Y(_0921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4081_ (.Y(_0922_),
    .A(_0919_),
    .B(_0920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4082_ (.Y(_0923_),
    .A(_0901_),
    .B(_0922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4083_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0874_),
    .A2(_0893_),
    .Y(_0924_),
    .B1(_0895_));
 sg13g2_or2_1 _4084_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0925_),
    .B(_0924_),
    .A(_0923_));
 sg13g2_xor2_1 _4085_ (.B(_0924_),
    .A(_0923_),
    .X(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4086_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0867_),
    .A2(_0898_),
    .Y(_0927_),
    .B1(_0897_));
 sg13g2_nor2b_1 _4087_ (.A(_0871_),
    .B_N(_0927_),
    .Y(_0928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4088_ (.B1(_0898_),
    .VDD(VPWR),
    .Y(_0929_),
    .VSS(VGND),
    .A1(_0868_),
    .A2(_0897_));
 sg13g2_a21oi_2 _4089_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0929_),
    .Y(_0930_),
    .A2(_0928_),
    .A1(_0870_));
 sg13g2_nand2_1 _4090_ (.Y(_0931_),
    .A(_0926_),
    .B(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4091_ (.B(_0930_),
    .A(_0926_),
    .X(_0119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4092_ (.A2(_0922_),
    .A1(_0901_),
    .B1(_0921_),
    .X(_0932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4093_ (.A2(_0914_),
    .A1(_0907_),
    .B1(_0916_),
    .X(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4094_ (.B1(_0911_),
    .VDD(VPWR),
    .Y(_0934_),
    .VSS(VGND),
    .A1(_0908_),
    .A2(_0912_));
 sg13g2_nand2_1 _4095_ (.Y(_0935_),
    .A(net966),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4096_ (.Y(_0936_),
    .A(net961),
    .B(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4097_ (.Y(_0937_),
    .A(net909),
    .B(net962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4098_ (.B(_0937_),
    .A(_0909_),
    .X(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4099_ (.Y(_0939_),
    .B(_0938_),
    .A_N(_0935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4100_ (.Y(_0940_),
    .A(_0935_),
    .B(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4101_ (.A(_0904_),
    .B_N(_0940_),
    .Y(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4102_ (.Y(_0942_),
    .A(_0904_),
    .B(_0940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4103_ (.Y(_0943_),
    .A(_0934_),
    .B(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4104_ (.A(_0903_),
    .B(_0943_),
    .Y(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4105_ (.B(_0943_),
    .A(_0903_),
    .X(_0945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4106_ (.Y(_0946_),
    .B(_0945_),
    .A_N(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4107_ (.Y(_0947_),
    .A(_0918_),
    .B(_0945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4108_ (.Y(_0948_),
    .A(_0933_),
    .B(_0947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4109_ (.B(_0947_),
    .A(_0933_),
    .X(_0949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4110_ (.Y(_0950_),
    .A(_0932_),
    .B(_0949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4111_ (.A(_0932_),
    .B(_0949_),
    .Y(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4112_ (.B(_0949_),
    .A(_0932_),
    .X(_0952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4113_ (.Y(_0953_),
    .A(_0925_),
    .B(_0931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4114_ (.B(_0953_),
    .A(_0952_),
    .X(_0120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4115_ (.A(_0926_),
    .B(_0952_),
    .X(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0925_),
    .A2(_0950_),
    .Y(_0955_),
    .B1(_0951_));
 sg13g2_a21o_1 _4117_ (.A2(_0954_),
    .A1(_0930_),
    .B1(_0955_),
    .X(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4118_ (.A(_0946_),
    .B(_0948_),
    .X(_0957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4119_ (.A2(_0942_),
    .A1(_0934_),
    .B1(_0941_),
    .X(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4120_ (.Y(_0959_),
    .A(net964),
    .B(\DP_2.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4121_ (.Y(_0960_),
    .A(net907),
    .B(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4122_ (.Y(_0961_),
    .A(net909),
    .B(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4123_ (.B(_0961_),
    .A(_0936_),
    .X(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4124_ (.Y(_0963_),
    .B(_0962_),
    .A_N(_0959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4125_ (.Y(_0964_),
    .A(_0959_),
    .B(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4126_ (.B1(_0939_),
    .VDD(VPWR),
    .Y(_0965_),
    .VSS(VGND),
    .A1(_0909_),
    .A2(_0937_));
 sg13g2_nand2_1 _4127_ (.Y(_0966_),
    .A(_0964_),
    .B(_0965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4128_ (.B(_0965_),
    .A(_0964_),
    .X(_0967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4129_ (.Y(_0968_),
    .A(_0944_),
    .B(_0967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4130_ (.A(_0968_),
    .B_N(_0958_),
    .Y(_0969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4131_ (.B(_0968_),
    .A(_0958_),
    .X(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4132_ (.A(_0957_),
    .B(_0970_),
    .Y(_0971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4133_ (.B(_0970_),
    .A(_0957_),
    .X(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4134_ (.B(_0972_),
    .A(_0956_),
    .X(_0121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4135_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0956_),
    .A2(_0972_),
    .Y(_0973_),
    .B1(_0971_));
 sg13g2_a21oi_1 _4136_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0944_),
    .A2(_0967_),
    .Y(_0974_),
    .B1(_0969_));
 sg13g2_o21ai_1 _4137_ (.B1(_0963_),
    .VDD(VPWR),
    .Y(_0975_),
    .VSS(VGND),
    .A1(_0936_),
    .A2(_0961_));
 sg13g2_nand2_1 _4138_ (.Y(_0976_),
    .A(net961),
    .B(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4139_ (.Y(_0977_),
    .A(_0960_),
    .B(_0976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4140_ (.Y(_0978_),
    .A(_0975_),
    .B(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4141_ (.Y(_0979_),
    .A(_0966_),
    .B(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4142_ (.Y(_0980_),
    .A(_0974_),
    .B(_0979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4143_ (.Y(_0122_),
    .A(_0973_),
    .B(_0980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4144_ (.A(net871),
    .B(net819),
    .X(_0079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4145_ (.X(_0981_),
    .A(net869),
    .B(net813),
    .C(_0079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4146_ (.Y(_0982_),
    .B1(net813),
    .B2(net871),
    .A2(net869),
    .A1(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4147_ (.A(_0981_),
    .B(_0982_),
    .Y(_0080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4148_ (.A(net871),
    .B(net811),
    .X(_0983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4149_ (.A(net819),
    .B(net869),
    .C(net813),
    .D(net867),
    .X(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4150_ (.Y(_0985_),
    .B1(net867),
    .B2(net819),
    .A2(net440),
    .A1(net869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4151_ (.A(_0984_),
    .B(_0985_),
    .Y(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4152_ (.B(_0986_),
    .A(_0983_),
    .X(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4153_ (.Y(_0988_),
    .A(_0981_),
    .B(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4154_ (.B(_0987_),
    .A(_0981_),
    .X(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4155_ (.Y(_0989_),
    .A(net363),
    .B(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4156_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0983_),
    .A2(_0986_),
    .Y(_0990_),
    .B1(_0984_));
 sg13g2_nand2_1 _4157_ (.Y(_0991_),
    .A(net869),
    .B(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4158_ (.A(net819),
    .B(net813),
    .C(net867),
    .D(net865),
    .X(_0992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4159_ (.B(net813),
    .C(net867),
    .A(net818),
    .Y(_0993_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net865));
 sg13g2_a22oi_1 _4160_ (.Y(_0994_),
    .B1(net865),
    .B2(net819),
    .A2(net867),
    .A1(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4161_ (.A(_0991_),
    .B(_0992_),
    .C(_0994_),
    .Y(_0995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4162_ (.B1(_0991_),
    .VDD(VPWR),
    .Y(_0996_),
    .VSS(VGND),
    .A1(_0992_),
    .A2(_0994_));
 sg13g2_nor2b_1 _4163_ (.A(_0995_),
    .B_N(_0996_),
    .Y(_0997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4164_ (.Y(_0998_),
    .B(_0997_),
    .A_N(_0990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4165_ (.Y(_0999_),
    .A(_0990_),
    .B(_0997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4166_ (.Y(_1000_),
    .B(_0999_),
    .A_N(_0989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4167_ (.Y(_1001_),
    .A(_0989_),
    .B(_0999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4168_ (.A(_0988_),
    .B_N(_1001_),
    .Y(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4169_ (.Y(_0082_),
    .A(_0988_),
    .B(_1001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4170_ (.Y(_1003_),
    .B1(net808),
    .B2(\DP_3.matrix[36] ),
    .A2(net809),
    .A1(net870),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4171_ (.Y(_1004_),
    .A(net870),
    .B(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4172_ (.A(_0989_),
    .B(_1004_),
    .Y(_1005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4173_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1006_),
    .B(_1005_),
    .A(_1003_));
 sg13g2_o21ai_1 _4174_ (.B1(_0993_),
    .VDD(VPWR),
    .Y(_1007_),
    .VSS(VGND),
    .A1(_0991_),
    .A2(_0994_));
 sg13g2_nand2_1 _4175_ (.Y(_1008_),
    .A(net867),
    .B(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4176_ (.A(net818),
    .B(net816),
    .C(net865),
    .D(net863),
    .X(_1009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4177_ (.B(net816),
    .C(net865),
    .A(net818),
    .Y(_1010_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net863));
 sg13g2_a22oi_1 _4178_ (.Y(_1011_),
    .B1(net863),
    .B2(net818),
    .A2(net865),
    .A1(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4179_ (.A(_1008_),
    .B(_1009_),
    .C(_1011_),
    .X(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4180_ (.B1(_1008_),
    .VDD(VPWR),
    .Y(_1013_),
    .VSS(VGND),
    .A1(_1009_),
    .A2(_1011_));
 sg13g2_nand3_1 _4181_ (.B(_1012_),
    .C(_1013_),
    .A(_1007_),
    .Y(_1014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4182_ (.A2(_1013_),
    .A1(_1012_),
    .B1(_1007_),
    .X(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4183_ (.Y(_1016_),
    .A(_1014_),
    .B(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4184_ (.B(_1016_),
    .A(_1006_),
    .X(_1017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4185_ (.Y(_1018_),
    .A(_0998_),
    .B(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4186_ (.Y(_1019_),
    .A(_1017_),
    .B(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4187_ (.B(_1018_),
    .A(_1017_),
    .X(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4188_ (.A(_1002_),
    .B(_1020_),
    .X(_1021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4189_ (.B(_1020_),
    .A(_1002_),
    .X(_0083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4190_ (.B1(_1014_),
    .VDD(VPWR),
    .Y(_1022_),
    .VSS(VGND),
    .A1(_1006_),
    .A2(_1016_));
 sg13g2_nand2_1 _4191_ (.Y(_1023_),
    .A(net871),
    .B(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4192_ (.Y(_1024_),
    .A(net868),
    .B(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4193_ (.Y(_1025_),
    .A(net868),
    .B(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4194_ (.B(_1025_),
    .A(_1004_),
    .X(_1026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4195_ (.Y(_1027_),
    .B(_1026_),
    .A_N(_1023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4196_ (.B(_1026_),
    .A(_1023_),
    .X(_1028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4197_ (.B1(_1010_),
    .VDD(VPWR),
    .Y(_1029_),
    .VSS(VGND),
    .A1(_1008_),
    .A2(_1011_));
 sg13g2_nand2_1 _4198_ (.Y(_1030_),
    .A(net812),
    .B(net866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4199_ (.A(net818),
    .B(net816),
    .C(net863),
    .D(net862),
    .X(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4200_ (.B(net816),
    .C(net863),
    .A(net818),
    .Y(_1032_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net862));
 sg13g2_a22oi_1 _4201_ (.Y(_1033_),
    .B1(net862),
    .B2(net818),
    .A2(net863),
    .A1(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4202_ (.A(_1030_),
    .B(_1031_),
    .C(_1033_),
    .X(_1034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4203_ (.B1(_1030_),
    .VDD(VPWR),
    .Y(_1035_),
    .VSS(VGND),
    .A1(_1031_),
    .A2(_1033_));
 sg13g2_and3_1 _4204_ (.X(_1036_),
    .A(_1029_),
    .B(_1034_),
    .C(_1035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4205_ (.B(_1034_),
    .C(_1035_),
    .A(_1029_),
    .Y(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4206_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1034_),
    .A2(_1035_),
    .Y(_1038_),
    .B1(_1029_));
 sg13g2_or3_1 _4207_ (.A(_1028_),
    .B(_1036_),
    .C(_1038_),
    .X(_1039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4208_ (.B1(_1028_),
    .VDD(VPWR),
    .Y(_1040_),
    .VSS(VGND),
    .A1(_1036_),
    .A2(_1038_));
 sg13g2_nand3_1 _4209_ (.B(_1039_),
    .C(_1040_),
    .A(_1022_),
    .Y(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4210_ (.A2(_1040_),
    .A1(_1039_),
    .B1(_1022_),
    .X(_1042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4211_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1041_),
    .A2(_1042_),
    .Y(_1043_),
    .B1(_1005_));
 sg13g2_and3_1 _4212_ (.X(_1044_),
    .A(_1005_),
    .B(_1041_),
    .C(_1042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4213_ (.B(_1041_),
    .C(_1042_),
    .A(_1005_),
    .Y(_1045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4214_ (.A(_1019_),
    .B(_1043_),
    .C(_1044_),
    .Y(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4215_ (.B1(_1019_),
    .VDD(VPWR),
    .Y(_1047_),
    .VSS(VGND),
    .A1(_1043_),
    .A2(_1044_));
 sg13g2_nand2b_1 _4216_ (.Y(_1048_),
    .B(_1047_),
    .A_N(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4217_ (.Y(_0127_),
    .A(_1021_),
    .B(_1048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4218_ (.Y(_1049_),
    .A(_1041_),
    .B(_1045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4219_ (.B1(_1027_),
    .VDD(VPWR),
    .Y(_1050_),
    .VSS(VGND),
    .A1(_1004_),
    .A2(_1025_));
 sg13g2_nand2_1 _4220_ (.Y(_1051_),
    .A(net871),
    .B(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4221_ (.Y(_1052_),
    .B(_1050_),
    .A_N(_1051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4222_ (.B(_1051_),
    .A(_1050_),
    .X(_1053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4223_ (.B1(_1037_),
    .VDD(VPWR),
    .Y(_1054_),
    .VSS(VGND),
    .A1(_1028_),
    .A2(_1038_));
 sg13g2_nand2_1 _4224_ (.Y(_1055_),
    .A(net870),
    .B(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4225_ (.Y(_1056_),
    .A(net866),
    .B(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4226_ (.Y(_1057_),
    .A(net866),
    .B(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4227_ (.B(_1057_),
    .A(_1024_),
    .X(_1058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4228_ (.Y(_1059_),
    .B(_1058_),
    .A_N(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4229_ (.Y(_1060_),
    .A(_1055_),
    .B(_1058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4230_ (.B1(_1032_),
    .VDD(VPWR),
    .Y(_1061_),
    .VSS(VGND),
    .A1(_1030_),
    .A2(_1033_));
 sg13g2_nand2_1 _4231_ (.Y(_1062_),
    .A(net812),
    .B(net864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4232_ (.A(net817),
    .B(net814),
    .C(net862),
    .D(net860),
    .X(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4233_ (.B(net814),
    .C(net862),
    .A(net817),
    .Y(_1064_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net860));
 sg13g2_a22oi_1 _4234_ (.Y(_1065_),
    .B1(net860),
    .B2(net817),
    .A2(net862),
    .A1(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4235_ (.A(_1062_),
    .B(_1063_),
    .C(_1065_),
    .X(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4236_ (.B1(_1062_),
    .VDD(VPWR),
    .Y(_1067_),
    .VSS(VGND),
    .A1(_1063_),
    .A2(_1065_));
 sg13g2_and3_1 _4237_ (.X(_1068_),
    .A(_1061_),
    .B(_1066_),
    .C(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4238_ (.B(_1066_),
    .C(_1067_),
    .A(_1061_),
    .Y(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4239_ (.A2(_1067_),
    .A1(_1066_),
    .B1(_1061_),
    .X(_1070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4240_ (.B(_1069_),
    .C(_1070_),
    .A(_1060_),
    .Y(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4241_ (.A2(_1070_),
    .A1(_1069_),
    .B1(_1060_),
    .X(_1072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4242_ (.B(_1071_),
    .C(_1072_),
    .A(_1054_),
    .Y(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4243_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1071_),
    .A2(_1072_),
    .Y(_1074_),
    .B1(_1054_));
 sg13g2_a21o_1 _4244_ (.A2(_1072_),
    .A1(_1071_),
    .B1(_1054_),
    .X(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4245_ (.Y(_1076_),
    .A(_1073_),
    .B(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4246_ (.Y(_1077_),
    .A(_1053_),
    .B(_1076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4247_ (.Y(_1078_),
    .B(_1049_),
    .A_N(_1077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4248_ (.B(_1077_),
    .A(_1049_),
    .X(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4249_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1021_),
    .A2(_1047_),
    .Y(_1080_),
    .B1(_1046_));
 sg13g2_xor2_1 _4250_ (.B(_1080_),
    .A(_1079_),
    .X(_0134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4251_ (.B1(_1073_),
    .VDD(VPWR),
    .Y(_1081_),
    .VSS(VGND),
    .A1(_1053_),
    .A2(_1074_));
 sg13g2_o21ai_1 _4252_ (.B1(_1059_),
    .VDD(VPWR),
    .Y(_1082_),
    .VSS(VGND),
    .A1(_1024_),
    .A2(_1057_));
 sg13g2_a22oi_1 _4253_ (.Y(_1083_),
    .B1(net801),
    .B2(\DP_3.matrix[36] ),
    .A2(net803),
    .A1(net869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4254_ (.Y(_1084_),
    .A(net870),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4255_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1085_),
    .B(_1084_),
    .A(_1051_));
 sg13g2_nor2b_1 _4256_ (.A(_1083_),
    .B_N(_1085_),
    .Y(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4257_ (.A(_1082_),
    .B(_1086_),
    .X(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4258_ (.Y(_1088_),
    .A(_1082_),
    .B(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4259_ (.A2(_1070_),
    .A1(_1060_),
    .B1(_1068_),
    .X(_1089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4260_ (.Y(_1090_),
    .A(net868),
    .B(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4261_ (.Y(_1091_),
    .A(net810),
    .B(net864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4262_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1092_),
    .B(_1091_),
    .A(_1056_));
 sg13g2_xnor2_1 _4263_ (.Y(_1093_),
    .A(_1056_),
    .B(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4264_ (.Y(_1094_),
    .A(_1090_),
    .B(_1093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4265_ (.B1(_1064_),
    .VDD(VPWR),
    .Y(_1095_),
    .VSS(VGND),
    .A1(_1062_),
    .A2(_1065_));
 sg13g2_nand2_1 _4266_ (.Y(_1096_),
    .A(net812),
    .B(net861),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4267_ (.A(net817),
    .B(net814),
    .C(net858),
    .D(net857),
    .X(_1097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4268_ (.B(net814),
    .C(net858),
    .A(net817),
    .Y(_1098_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net855));
 sg13g2_a22oi_1 _4269_ (.Y(_1099_),
    .B1(net855),
    .B2(\DP_4.matrix[36] ),
    .A2(net858),
    .A1(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4270_ (.A(_1096_),
    .B(_1097_),
    .C(_1099_),
    .X(_1100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4271_ (.B1(_1096_),
    .VDD(VPWR),
    .Y(_1101_),
    .VSS(VGND),
    .A1(_1097_),
    .A2(_1099_));
 sg13g2_and3_1 _4272_ (.X(_1102_),
    .A(_1095_),
    .B(_1100_),
    .C(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4273_ (.B(_1100_),
    .C(_1101_),
    .A(_1095_),
    .Y(_1103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4274_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1100_),
    .A2(_1101_),
    .Y(_1104_),
    .B1(_1095_));
 sg13g2_or3_1 _4275_ (.A(_1094_),
    .B(_1102_),
    .C(_1104_),
    .X(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4276_ (.B1(_1094_),
    .VDD(VPWR),
    .Y(_1106_),
    .VSS(VGND),
    .A1(_1102_),
    .A2(_1104_));
 sg13g2_and3_1 _4277_ (.X(_1107_),
    .A(_1089_),
    .B(_1105_),
    .C(_1106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4278_ (.B(_1105_),
    .C(_1106_),
    .A(_1089_),
    .Y(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4279_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1105_),
    .A2(_1106_),
    .Y(_1109_),
    .B1(_1089_));
 sg13g2_or3_1 _4280_ (.A(_1088_),
    .B(_1107_),
    .C(_1109_),
    .X(_1110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4281_ (.B1(_1088_),
    .VDD(VPWR),
    .Y(_1111_),
    .VSS(VGND),
    .A1(_1107_),
    .A2(_1109_));
 sg13g2_nand3_1 _4282_ (.B(_1110_),
    .C(_1111_),
    .A(_1081_),
    .Y(_1112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4283_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1110_),
    .A2(_1111_),
    .Y(_1113_),
    .B1(_1081_));
 sg13g2_a21o_1 _4284_ (.A2(_1111_),
    .A1(_1110_),
    .B1(_1081_),
    .X(_1114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4285_ (.Y(_1115_),
    .A(_1112_),
    .B(_1114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4286_ (.B(_1115_),
    .A(_1052_),
    .X(_1116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4287_ (.B1(_1078_),
    .VDD(VPWR),
    .Y(_1117_),
    .VSS(VGND),
    .A1(_1079_),
    .A2(_1080_));
 sg13g2_nand2_1 _4288_ (.Y(_1118_),
    .A(_1116_),
    .B(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4289_ (.B(_1117_),
    .A(_1116_),
    .X(_0135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4290_ (.B1(_1108_),
    .VDD(VPWR),
    .Y(_1119_),
    .VSS(VGND),
    .A1(_1088_),
    .A2(_1109_));
 sg13g2_o21ai_1 _4291_ (.B1(_1092_),
    .VDD(VPWR),
    .Y(_1120_),
    .VSS(VGND),
    .A1(_1090_),
    .A2(_1093_));
 sg13g2_nand2_1 _4292_ (.Y(_1121_),
    .A(net871),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4293_ (.Y(_1122_),
    .A(net868),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4294_ (.Y(_1123_),
    .A(net868),
    .B(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4295_ (.B(_1123_),
    .A(_1084_),
    .X(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4296_ (.Y(_1125_),
    .B(_1124_),
    .A_N(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4297_ (.Y(_1126_),
    .A(_1121_),
    .B(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4298_ (.Y(_1127_),
    .A(_1120_),
    .B(_1126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4299_ (.Y(_1128_),
    .A(_1120_),
    .B(_1126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4300_ (.Y(_1129_),
    .A(_1085_),
    .B(_1128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4301_ (.B1(_1103_),
    .VDD(VPWR),
    .Y(_1130_),
    .VSS(VGND),
    .A1(_1094_),
    .A2(_1104_));
 sg13g2_nand2_1 _4302_ (.Y(_1131_),
    .A(net866),
    .B(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4303_ (.Y(_1132_),
    .A(net807),
    .B(net861),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4304_ (.A(net809),
    .B(\DP_3.matrix[40] ),
    .C(net807),
    .D(\DP_3.matrix[41] ),
    .X(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4305_ (.Y(_1134_),
    .B1(net861),
    .B2(net809),
    .A2(net808),
    .A1(net864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4306_ (.A(_1131_),
    .B(_1133_),
    .C(_1134_),
    .Y(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4307_ (.B1(_1131_),
    .VDD(VPWR),
    .Y(_1136_),
    .VSS(VGND),
    .A1(_1133_),
    .A2(_1134_));
 sg13g2_nand2b_1 _4308_ (.Y(_1137_),
    .B(_1136_),
    .A_N(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4309_ (.B1(_1098_),
    .VDD(VPWR),
    .Y(_1138_),
    .VSS(VGND),
    .A1(_1096_),
    .A2(_1099_));
 sg13g2_nand2_1 _4310_ (.Y(_1139_),
    .A(net811),
    .B(net858),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4311_ (.A(net817),
    .B(net814),
    .C(net855),
    .D(net999),
    .X(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4312_ (.B(net814),
    .C(net855),
    .A(net817),
    .Y(_1141_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net999));
 sg13g2_a22oi_1 _4313_ (.Y(_1142_),
    .B1(net999),
    .B2(net817),
    .A2(net855),
    .A1(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4314_ (.A(_1139_),
    .B(_1140_),
    .C(_1142_),
    .X(_1143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4315_ (.B1(_1139_),
    .VDD(VPWR),
    .Y(_1144_),
    .VSS(VGND),
    .A1(_1140_),
    .A2(_1142_));
 sg13g2_and3_1 _4316_ (.X(_1145_),
    .A(_1138_),
    .B(_1143_),
    .C(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4317_ (.B(_1143_),
    .C(_1144_),
    .A(_1138_),
    .Y(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4318_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1143_),
    .A2(_1144_),
    .Y(_1147_),
    .B1(_1138_));
 sg13g2_or3_1 _4319_ (.A(_1137_),
    .B(_1145_),
    .C(_1147_),
    .X(_1148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4320_ (.B1(_1137_),
    .VDD(VPWR),
    .Y(_1149_),
    .VSS(VGND),
    .A1(_1145_),
    .A2(_1147_));
 sg13g2_and3_1 _4321_ (.X(_1150_),
    .A(_1130_),
    .B(_1148_),
    .C(_1149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4322_ (.B(_1148_),
    .C(_1149_),
    .A(_1130_),
    .Y(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4323_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1148_),
    .A2(_1149_),
    .Y(_1152_),
    .B1(_1130_));
 sg13g2_or3_1 _4324_ (.A(_1129_),
    .B(_1150_),
    .C(_1152_),
    .X(_1153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4325_ (.B1(_1129_),
    .VDD(VPWR),
    .Y(_1154_),
    .VSS(VGND),
    .A1(_1150_),
    .A2(_1152_));
 sg13g2_nand3_1 _4326_ (.B(_1153_),
    .C(_1154_),
    .A(_1119_),
    .Y(_1155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4327_ (.A2(_1154_),
    .A1(_1153_),
    .B1(_1119_),
    .X(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4328_ (.A2(_1156_),
    .A1(_1155_),
    .B1(_1087_),
    .X(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4329_ (.B(_1155_),
    .C(_1156_),
    .A(_1087_),
    .Y(_1158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4330_ (.B1(_1112_),
    .VDD(VPWR),
    .Y(_1159_),
    .VSS(VGND),
    .A1(_1052_),
    .A2(_1113_));
 sg13g2_nand3_1 _4331_ (.B(_1158_),
    .C(_1159_),
    .A(_1157_),
    .Y(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4332_ (.A2(_1158_),
    .A1(_1157_),
    .B1(_1159_),
    .X(_1161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4333_ (.A(_1160_),
    .B(_1161_),
    .X(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4334_ (.B(_1117_),
    .C(_1162_),
    .A(_1116_),
    .Y(_1163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4335_ (.Y(_0136_),
    .A(_1118_),
    .B(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4336_ (.B1(_1127_),
    .VDD(VPWR),
    .Y(_1164_),
    .VSS(VGND),
    .A1(_1085_),
    .A2(_1128_));
 sg13g2_o21ai_1 _4337_ (.B1(_1151_),
    .VDD(VPWR),
    .Y(_1165_),
    .VSS(VGND),
    .A1(_1129_),
    .A2(_1152_));
 sg13g2_o21ai_1 _4338_ (.B1(_1125_),
    .VDD(VPWR),
    .Y(_1166_),
    .VSS(VGND),
    .A1(_1084_),
    .A2(_1123_));
 sg13g2_or2_1 _4339_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1167_),
    .B(_1135_),
    .A(_1133_));
 sg13g2_nand2_1 _4340_ (.Y(_1168_),
    .A(net870),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4341_ (.Y(_1169_),
    .A(net866),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4342_ (.Y(_1170_),
    .A(net866),
    .B(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4343_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1171_),
    .B(_1169_),
    .A(_1123_));
 sg13g2_xnor2_1 _4344_ (.Y(_1172_),
    .A(_1122_),
    .B(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4345_ (.B(_1172_),
    .A(_1168_),
    .X(_1173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4346_ (.Y(_1174_),
    .A(_1167_),
    .B(_1173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4347_ (.A(_1174_),
    .B_N(_1166_),
    .Y(_1175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4348_ (.B(_1174_),
    .A(_1166_),
    .X(_1176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4349_ (.B1(_1146_),
    .VDD(VPWR),
    .Y(_1177_),
    .VSS(VGND),
    .A1(_1137_),
    .A2(_1147_));
 sg13g2_nand2_1 _4350_ (.Y(_1178_),
    .A(net864),
    .B(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4351_ (.Y(_1179_),
    .A(net809),
    .B(net858),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4352_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1180_),
    .B(_1179_),
    .A(_1132_));
 sg13g2_and2_1 _4353_ (.A(_1132_),
    .B(_1179_),
    .X(_1181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4354_ (.Y(_1182_),
    .A(_1132_),
    .B(_1179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4355_ (.Y(_1183_),
    .A(_1178_),
    .B(_1182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4356_ (.B1(_1141_),
    .VDD(VPWR),
    .Y(_1184_),
    .VSS(VGND),
    .A1(_1139_),
    .A2(_1142_));
 sg13g2_nand2_1 _4357_ (.Y(_1185_),
    .A(net812),
    .B(net999),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4358_ (.A(net815),
    .B(net811),
    .C(net855),
    .D(net999),
    .X(_1186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4359_ (.Y(_1187_),
    .B1(net999),
    .B2(net815),
    .A2(net855),
    .A1(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4360_ (.A(_1186_),
    .B(_1187_),
    .Y(_1188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4361_ (.Y(_1189_),
    .A(_1184_),
    .B(_1188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4362_ (.Y(_1190_),
    .A(_1184_),
    .B(_1188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4363_ (.B(_1190_),
    .A(_1183_),
    .X(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4364_ (.Y(_1192_),
    .A(_1177_),
    .B(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4365_ (.Y(_1193_),
    .A(_1177_),
    .B(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4366_ (.B(_1193_),
    .A(_1176_),
    .X(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4367_ (.Y(_1195_),
    .A(_1165_),
    .B(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4368_ (.Y(_1196_),
    .A(_1165_),
    .B(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4369_ (.Y(_1197_),
    .B(_1164_),
    .A_N(_1196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4370_ (.B(_1196_),
    .A(_1164_),
    .X(_1198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4371_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1155_),
    .A2(_1158_),
    .Y(_1199_),
    .B1(_1198_));
 sg13g2_a21o_1 _4372_ (.A2(_1158_),
    .A1(_1155_),
    .B1(_1198_),
    .X(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4373_ (.X(_1201_),
    .A(_1155_),
    .B(_1158_),
    .C(_1198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4374_ (.A(_1199_),
    .B(_1201_),
    .Y(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4375_ (.Y(_1203_),
    .A(_1160_),
    .B(_1163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4376_ (.B(_1203_),
    .A(_1202_),
    .X(_0137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4377_ (.A2(_1173_),
    .A1(_1167_),
    .B1(_1175_),
    .X(_1204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4378_ (.B1(_1192_),
    .VDD(VPWR),
    .Y(_1205_),
    .VSS(VGND),
    .A1(_1176_),
    .A2(_1193_));
 sg13g2_o21ai_1 _4379_ (.B1(_1171_),
    .VDD(VPWR),
    .Y(_1206_),
    .VSS(VGND),
    .A1(_1168_),
    .A2(_1172_));
 sg13g2_o21ai_1 _4380_ (.B1(_1180_),
    .VDD(VPWR),
    .Y(_1207_),
    .VSS(VGND),
    .A1(_1178_),
    .A2(_1181_));
 sg13g2_nand2_1 _4381_ (.Y(_1208_),
    .A(net868),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4382_ (.Y(_1209_),
    .A(net864),
    .B(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4383_ (.Y(_1210_),
    .A(net864),
    .B(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4384_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1211_),
    .B(_1209_),
    .A(_1170_));
 sg13g2_xnor2_1 _4385_ (.Y(_1212_),
    .A(_1169_),
    .B(_1210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4386_ (.B(_1212_),
    .A(_1208_),
    .X(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4387_ (.Y(_1214_),
    .A(_1207_),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4388_ (.A(_1214_),
    .B_N(_1206_),
    .Y(_1215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4389_ (.B(_1214_),
    .A(_1206_),
    .X(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4390_ (.B1(_1189_),
    .VDD(VPWR),
    .Y(_1217_),
    .VSS(VGND),
    .A1(_1183_),
    .A2(_1190_));
 sg13g2_a21oi_1 _4391_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net815),
    .A2(net855),
    .Y(_1218_),
    .B1(_1185_));
 sg13g2_nand2_1 _4392_ (.Y(_1219_),
    .A(net861),
    .B(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4393_ (.Y(_1220_),
    .A(net807),
    .B(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4394_ (.A(net810),
    .B(net807),
    .C(net859),
    .D(net856),
    .X(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4395_ (.Y(_1222_),
    .B1(net856),
    .B2(net810),
    .A2(net859),
    .A1(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4396_ (.A(_1219_),
    .B(_1221_),
    .C(_1222_),
    .Y(_1223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4397_ (.B1(_1219_),
    .VDD(VPWR),
    .Y(_1224_),
    .VSS(VGND),
    .A1(_1221_),
    .A2(_1222_));
 sg13g2_nor2b_1 _4398_ (.A(_1223_),
    .B_N(_1224_),
    .Y(_1225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4399_ (.Y(_1226_),
    .A(_1218_),
    .B(_1225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4400_ (.Y(_1227_),
    .B(_1217_),
    .A_N(_1226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4401_ (.B(_1226_),
    .A(_1217_),
    .X(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4402_ (.B(_1228_),
    .A(_1216_),
    .X(_1229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4403_ (.Y(_1230_),
    .A(_1205_),
    .B(_1229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4404_ (.B(_1229_),
    .A(_1205_),
    .X(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4405_ (.Y(_1232_),
    .A(_1204_),
    .B(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4406_ (.Y(_1233_),
    .A(_1204_),
    .B(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4407_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1195_),
    .A2(_1197_),
    .Y(_1234_),
    .B1(_1233_));
 sg13g2_nand3_1 _4408_ (.B(_1197_),
    .C(_1233_),
    .A(_1195_),
    .Y(_1235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4409_ (.A(_1234_),
    .B_N(_1235_),
    .Y(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4410_ (.B(_1117_),
    .C(_1162_),
    .A(_1116_),
    .Y(_1237_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1202_));
 sg13g2_a21oi_1 _4411_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1160_),
    .A2(_1200_),
    .Y(_1238_),
    .B1(_1201_));
 sg13g2_nand2b_1 _4412_ (.Y(_1239_),
    .B(_1237_),
    .A_N(_1238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4413_ (.B(_1239_),
    .A(_1236_),
    .X(_0128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4414_ (.A2(_1213_),
    .A1(_1207_),
    .B1(_1215_),
    .X(_1240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4415_ (.B1(_1227_),
    .VDD(VPWR),
    .Y(_1241_),
    .VSS(VGND),
    .A1(_1216_),
    .A2(_1228_));
 sg13g2_a21o_1 _4416_ (.A2(_1225_),
    .A1(_1218_),
    .B1(_1186_),
    .X(_1242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4417_ (.Y(_1243_),
    .A(net805),
    .B(net859),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4418_ (.Y(_1244_),
    .A(net810),
    .B(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4419_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1245_),
    .B(_1244_),
    .A(_1220_));
 sg13g2_xnor2_1 _4420_ (.Y(_1246_),
    .A(_1220_),
    .B(_1244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4421_ (.B(_1246_),
    .A(_1243_),
    .X(_1247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4422_ (.Y(_1248_),
    .A(_1242_),
    .B(_1247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4423_ (.B1(_1211_),
    .VDD(VPWR),
    .Y(_1249_),
    .VSS(VGND),
    .A1(_1208_),
    .A2(_1212_));
 sg13g2_or2_1 _4424_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1250_),
    .B(_1223_),
    .A(_1221_));
 sg13g2_nand2_1 _4425_ (.Y(_1251_),
    .A(net866),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4426_ (.Y(_1252_),
    .A(net861),
    .B(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4427_ (.Y(_1253_),
    .A(net861),
    .B(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4428_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1254_),
    .B(_1252_),
    .A(_1210_));
 sg13g2_xnor2_1 _4429_ (.Y(_1255_),
    .A(_1209_),
    .B(_1253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4430_ (.B(_1255_),
    .A(_1251_),
    .X(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4431_ (.Y(_1257_),
    .A(_1250_),
    .B(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4432_ (.A(_1257_),
    .B_N(_1249_),
    .Y(_1258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4433_ (.B(_1257_),
    .A(_1249_),
    .X(_1259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4434_ (.A(_1248_),
    .B(_1259_),
    .Y(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4435_ (.B(_1259_),
    .A(_1248_),
    .X(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4436_ (.Y(_1262_),
    .A(_1241_),
    .B(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4437_ (.A(_1262_),
    .B_N(_1240_),
    .Y(_1263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4438_ (.B(_1262_),
    .A(_1240_),
    .X(_1264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1230_),
    .A2(_1232_),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_nand3_1 _4440_ (.B(_1232_),
    .C(_1264_),
    .A(_1230_),
    .Y(_1266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4441_ (.A(_1265_),
    .B_N(_1266_),
    .Y(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4442_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1236_),
    .A2(_1239_),
    .Y(_1268_),
    .B1(_1234_));
 sg13g2_xnor2_1 _4443_ (.Y(_0129_),
    .A(_1267_),
    .B(_1268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4444_ (.A2(_1256_),
    .A1(_1250_),
    .B1(_1258_),
    .X(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4445_ (.Y(_1270_),
    .B1(net1000),
    .B2(net807),
    .A2(net856),
    .A1(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4446_ (.Y(_1271_),
    .A(net805),
    .B(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4447_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1272_),
    .B(_1271_),
    .A(_1220_));
 sg13g2_nand2b_1 _4448_ (.Y(_1273_),
    .B(_1272_),
    .A_N(_1270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4449_ (.B1(_1254_),
    .VDD(VPWR),
    .Y(_1274_),
    .VSS(VGND),
    .A1(_1251_),
    .A2(_1255_));
 sg13g2_o21ai_1 _4450_ (.B1(_1245_),
    .VDD(VPWR),
    .Y(_1275_),
    .VSS(VGND),
    .A1(_1243_),
    .A2(_1246_));
 sg13g2_nand2_1 _4451_ (.Y(_1276_),
    .A(net864),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4452_ (.Y(_1277_),
    .A(net858),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4453_ (.Y(_1278_),
    .A(net859),
    .B(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4454_ (.B(_1278_),
    .A(_1252_),
    .X(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4455_ (.Y(_1280_),
    .B(_1279_),
    .A_N(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4456_ (.Y(_1281_),
    .A(_1276_),
    .B(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4457_ (.Y(_1282_),
    .A(_1275_),
    .B(_1281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4458_ (.A(_1282_),
    .B_N(_1274_),
    .Y(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4459_ (.B(_1282_),
    .A(_1274_),
    .X(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4460_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1285_),
    .B(_1284_),
    .A(_1273_));
 sg13g2_xor2_1 _4461_ (.B(_1284_),
    .A(_1273_),
    .X(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4462_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1242_),
    .A2(_1247_),
    .Y(_1287_),
    .B1(_1260_));
 sg13g2_nor2b_1 _4463_ (.A(_1287_),
    .B_N(_1286_),
    .Y(_1288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4464_ (.Y(_1289_),
    .A(_1286_),
    .B(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4465_ (.Y(_1290_),
    .A(_1269_),
    .B(_1289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4466_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1241_),
    .A2(_1261_),
    .Y(_1291_),
    .B1(_1263_));
 sg13g2_or2_1 _4467_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1292_),
    .B(_1291_),
    .A(_1290_));
 sg13g2_xor2_1 _4468_ (.B(_1291_),
    .A(_1290_),
    .X(_1293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4469_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1234_),
    .A2(_1266_),
    .Y(_1294_),
    .B1(_1265_));
 sg13g2_nor2b_1 _4470_ (.A(_1238_),
    .B_N(_1294_),
    .Y(_1295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4471_ (.B1(_1266_),
    .VDD(VPWR),
    .Y(_1296_),
    .VSS(VGND),
    .A1(_1235_),
    .A2(_1265_));
 sg13g2_a21oi_2 _4472_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1296_),
    .Y(_1297_),
    .A2(_1295_),
    .A1(_1237_));
 sg13g2_nand2_1 _4473_ (.Y(_1298_),
    .A(_1293_),
    .B(_1297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4474_ (.B(_1297_),
    .A(_1293_),
    .X(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4475_ (.A2(_1289_),
    .A1(_1269_),
    .B1(_1288_),
    .X(_1299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4476_ (.A2(_1281_),
    .A1(_1275_),
    .B1(_1283_),
    .X(_1300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4477_ (.B1(_1280_),
    .VDD(VPWR),
    .Y(_1301_),
    .VSS(VGND),
    .A1(_1252_),
    .A2(_1278_));
 sg13g2_nand2_1 _4478_ (.Y(_1302_),
    .A(net861),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4479_ (.Y(_1303_),
    .A(net856),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4480_ (.Y(_1304_),
    .A(net803),
    .B(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4481_ (.B(_1304_),
    .A(_1277_),
    .X(_1305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4482_ (.Y(_1306_),
    .B(_1305_),
    .A_N(_1302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4483_ (.Y(_1307_),
    .A(_1302_),
    .B(_1305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4484_ (.A(_1272_),
    .B_N(_1307_),
    .Y(_1308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4485_ (.Y(_1309_),
    .A(_1272_),
    .B(_1307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4486_ (.Y(_1310_),
    .A(_1301_),
    .B(_1309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4487_ (.A(_1271_),
    .B(_1310_),
    .Y(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4488_ (.B(_1310_),
    .A(_1271_),
    .X(_1312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4489_ (.Y(_1313_),
    .B(_1312_),
    .A_N(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4490_ (.Y(_1314_),
    .A(_1285_),
    .B(_1312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4491_ (.Y(_1315_),
    .A(_1300_),
    .B(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4492_ (.B(_1314_),
    .A(_1300_),
    .X(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4493_ (.Y(_1317_),
    .A(_1299_),
    .B(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4494_ (.A(_1299_),
    .B(_1316_),
    .Y(_1318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4495_ (.B(_1316_),
    .A(_1299_),
    .X(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4496_ (.Y(_1320_),
    .A(_1292_),
    .B(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4497_ (.B(_1320_),
    .A(_1319_),
    .X(_0131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4498_ (.A(_1293_),
    .B(_1319_),
    .X(_1321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4499_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1292_),
    .A2(_1317_),
    .Y(_1322_),
    .B1(_1318_));
 sg13g2_a21o_1 _4500_ (.A2(_1321_),
    .A1(_1297_),
    .B1(_1322_),
    .X(_1323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4501_ (.A(_1313_),
    .B(_1315_),
    .X(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4502_ (.A2(_1309_),
    .A1(_1301_),
    .B1(_1308_),
    .X(_1325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4503_ (.Y(_1326_),
    .A(net858),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4504_ (.Y(_1327_),
    .A(net801),
    .B(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4505_ (.Y(_1328_),
    .A(net803),
    .B(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4506_ (.B(_1328_),
    .A(_1303_),
    .X(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4507_ (.Y(_1330_),
    .B(_1329_),
    .A_N(_1326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4508_ (.Y(_1331_),
    .A(_1326_),
    .B(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4509_ (.B1(_1306_),
    .VDD(VPWR),
    .Y(_1332_),
    .VSS(VGND),
    .A1(_1277_),
    .A2(_1304_));
 sg13g2_nand2_1 _4510_ (.Y(_1333_),
    .A(_1331_),
    .B(_1332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4511_ (.B(_1332_),
    .A(_1331_),
    .X(_1334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4512_ (.Y(_1335_),
    .A(_1311_),
    .B(_1334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4513_ (.A(_1335_),
    .B_N(_1325_),
    .Y(_1336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4514_ (.B(_1335_),
    .A(_1325_),
    .X(_1337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4515_ (.A(_1324_),
    .B(_1337_),
    .Y(_1338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4516_ (.B(_1337_),
    .A(_1324_),
    .X(_1339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4517_ (.B(_1339_),
    .A(_1323_),
    .X(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1323_),
    .A2(_1339_),
    .Y(_1340_),
    .B1(_1338_));
 sg13g2_a21oi_1 _4519_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1311_),
    .A2(_1334_),
    .Y(_1341_),
    .B1(_1336_));
 sg13g2_o21ai_1 _4520_ (.B1(_1330_),
    .VDD(VPWR),
    .Y(_1342_),
    .VSS(VGND),
    .A1(_1304_),
    .A2(_1327_));
 sg13g2_nand2_1 _4521_ (.Y(_1343_),
    .A(net856),
    .B(\DP_4.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4522_ (.Y(_1344_),
    .A(_1327_),
    .B(_1343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4523_ (.Y(_1345_),
    .A(_1342_),
    .B(_1344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4524_ (.Y(_1346_),
    .A(_1333_),
    .B(_1345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4525_ (.Y(_1347_),
    .A(_1341_),
    .B(_1346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4526_ (.Y(_0133_),
    .A(_1340_),
    .B(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4527_ (.A(net886),
    .B(net833),
    .X(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4528_ (.X(_1348_),
    .A(net884),
    .B(net829),
    .C(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4529_ (.Y(_1349_),
    .B1(net829),
    .B2(net886),
    .A2(net884),
    .A1(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4530_ (.A(_1348_),
    .B(_1349_),
    .Y(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4531_ (.A(net886),
    .B(net827),
    .X(_1350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4532_ (.A(net833),
    .B(net884),
    .C(net829),
    .D(net882),
    .X(_1351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4533_ (.Y(_1352_),
    .B1(net882),
    .B2(net833),
    .A2(net829),
    .A1(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4534_ (.A(_1351_),
    .B(_1352_),
    .Y(_1353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4535_ (.B(_1353_),
    .A(_1350_),
    .X(_1354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4536_ (.Y(_1355_),
    .A(_1348_),
    .B(_1354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4537_ (.B(_1354_),
    .A(_1348_),
    .X(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4538_ (.Y(_1356_),
    .A(net886),
    .B(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4539_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1350_),
    .A2(_1353_),
    .Y(_1357_),
    .B1(_1351_));
 sg13g2_nand2_1 _4540_ (.Y(_1358_),
    .A(net884),
    .B(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4541_ (.A(net833),
    .B(net829),
    .C(net882),
    .D(net880),
    .X(_1359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4542_ (.B(net830),
    .C(net882),
    .A(net833),
    .Y(_1360_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net880));
 sg13g2_a22oi_1 _4543_ (.Y(_1361_),
    .B1(net880),
    .B2(net834),
    .A2(net882),
    .A1(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4544_ (.A(_1358_),
    .B(_1359_),
    .C(_1361_),
    .Y(_1362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4545_ (.B1(_1358_),
    .VDD(VPWR),
    .Y(_1363_),
    .VSS(VGND),
    .A1(_1359_),
    .A2(_1361_));
 sg13g2_nor2b_1 _4546_ (.A(_1362_),
    .B_N(_1363_),
    .Y(_1364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4547_ (.Y(_1365_),
    .B(_1364_),
    .A_N(_1357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4548_ (.Y(_1366_),
    .A(_1357_),
    .B(_1364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4549_ (.Y(_1367_),
    .B(_1366_),
    .A_N(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4550_ (.Y(_1368_),
    .A(_1356_),
    .B(_1366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4551_ (.A(_1355_),
    .B_N(_1368_),
    .Y(_1369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4552_ (.Y(_0087_),
    .A(_1355_),
    .B(_1368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4553_ (.Y(_1370_),
    .B1(net824),
    .B2(net886),
    .A2(net825),
    .A1(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4554_ (.Y(_1371_),
    .A(net885),
    .B(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4555_ (.A(_1356_),
    .B(_1371_),
    .Y(_1372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4556_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1373_),
    .B(_1372_),
    .A(_1370_));
 sg13g2_o21ai_1 _4557_ (.B1(_1360_),
    .VDD(VPWR),
    .Y(_1374_),
    .VSS(VGND),
    .A1(_1358_),
    .A2(_1361_));
 sg13g2_nand2_1 _4558_ (.Y(_1375_),
    .A(net883),
    .B(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4559_ (.A(net834),
    .B(net830),
    .C(net880),
    .D(net878),
    .X(_1376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4560_ (.B(net830),
    .C(net880),
    .A(net834),
    .Y(_1377_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net878));
 sg13g2_a22oi_1 _4561_ (.Y(_1378_),
    .B1(net878),
    .B2(net834),
    .A2(net880),
    .A1(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4562_ (.A(_1375_),
    .B(_1376_),
    .C(_1378_),
    .X(_1379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4563_ (.B1(_1375_),
    .VDD(VPWR),
    .Y(_1380_),
    .VSS(VGND),
    .A1(_1376_),
    .A2(_1378_));
 sg13g2_nand3_1 _4564_ (.B(_1379_),
    .C(_1380_),
    .A(_1374_),
    .Y(_1381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4565_ (.A2(_1380_),
    .A1(_1379_),
    .B1(_1374_),
    .X(_1382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4566_ (.Y(_1383_),
    .A(_1381_),
    .B(_1382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4567_ (.B(_1383_),
    .A(_1373_),
    .X(_1384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4568_ (.Y(_1385_),
    .A(_1365_),
    .B(_1367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4569_ (.Y(_1386_),
    .A(_1384_),
    .B(_1385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4570_ (.B(_1385_),
    .A(_1384_),
    .X(_1387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4571_ (.A(_1369_),
    .B(_1387_),
    .X(_1388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4572_ (.B(_1387_),
    .A(_1369_),
    .X(_0088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4573_ (.B1(_1381_),
    .VDD(VPWR),
    .Y(_1389_),
    .VSS(VGND),
    .A1(_1373_),
    .A2(_1383_));
 sg13g2_nand2_1 _4574_ (.Y(_1390_),
    .A(net886),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4575_ (.Y(_1391_),
    .A(net883),
    .B(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4576_ (.Y(_1392_),
    .A(net882),
    .B(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4577_ (.B(_1392_),
    .A(_1371_),
    .X(_1393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4578_ (.Y(_1394_),
    .B(_1393_),
    .A_N(_1390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4579_ (.B(_1393_),
    .A(_1390_),
    .X(_1395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4580_ (.B1(_1377_),
    .VDD(VPWR),
    .Y(_1396_),
    .VSS(VGND),
    .A1(_1375_),
    .A2(_1378_));
 sg13g2_nand2_1 _4581_ (.Y(_1397_),
    .A(net827),
    .B(net881),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4582_ (.A(net835),
    .B(net832),
    .C(net878),
    .D(net876),
    .X(_1398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4583_ (.B(net832),
    .C(net878),
    .A(net835),
    .Y(_1399_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net876));
 sg13g2_a22oi_1 _4584_ (.Y(_1400_),
    .B1(net876),
    .B2(net835),
    .A2(net879),
    .A1(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4585_ (.A(_1397_),
    .B(_1398_),
    .C(_1400_),
    .X(_1401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4586_ (.B1(_1397_),
    .VDD(VPWR),
    .Y(_1402_),
    .VSS(VGND),
    .A1(_1398_),
    .A2(_1400_));
 sg13g2_and3_1 _4587_ (.X(_1403_),
    .A(_1396_),
    .B(_1401_),
    .C(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4588_ (.B(_1401_),
    .C(_1402_),
    .A(_1396_),
    .Y(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4589_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1401_),
    .A2(_1402_),
    .Y(_1405_),
    .B1(_1396_));
 sg13g2_or3_1 _4590_ (.A(_1395_),
    .B(_1403_),
    .C(_1405_),
    .X(_1406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4591_ (.B1(_1395_),
    .VDD(VPWR),
    .Y(_1407_),
    .VSS(VGND),
    .A1(_1403_),
    .A2(_1405_));
 sg13g2_nand3_1 _4592_ (.B(_1406_),
    .C(_1407_),
    .A(_1389_),
    .Y(_1408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4593_ (.A2(_1407_),
    .A1(_1406_),
    .B1(_1389_),
    .X(_1409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4594_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1408_),
    .A2(_1409_),
    .Y(_1410_),
    .B1(_1372_));
 sg13g2_and3_1 _4595_ (.X(_1411_),
    .A(_1372_),
    .B(_1408_),
    .C(_1409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4596_ (.B(_1408_),
    .C(_1409_),
    .A(_1372_),
    .Y(_1412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4597_ (.A(_1386_),
    .B(_1410_),
    .C(_1411_),
    .Y(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4598_ (.B1(_1386_),
    .VDD(VPWR),
    .Y(_1414_),
    .VSS(VGND),
    .A1(_1410_),
    .A2(_1411_));
 sg13g2_nand2b_1 _4599_ (.Y(_1415_),
    .B(_1414_),
    .A_N(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4600_ (.Y(_0138_),
    .A(_1388_),
    .B(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4601_ (.Y(_1416_),
    .A(_1408_),
    .B(_1412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4602_ (.B1(_1394_),
    .VDD(VPWR),
    .Y(_1417_),
    .VSS(VGND),
    .A1(_1371_),
    .A2(_1392_));
 sg13g2_nand2_1 _4603_ (.Y(_1418_),
    .A(\DP_3.matrix[0] ),
    .B(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4604_ (.Y(_1419_),
    .B(_1417_),
    .A_N(_1418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4605_ (.B(_1418_),
    .A(_1417_),
    .X(_1420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4606_ (.B1(_1404_),
    .VDD(VPWR),
    .Y(_1421_),
    .VSS(VGND),
    .A1(_1395_),
    .A2(_1405_));
 sg13g2_nand2_1 _4607_ (.Y(_1422_),
    .A(net885),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4608_ (.Y(_1423_),
    .A(net881),
    .B(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4609_ (.Y(_1424_),
    .A(net881),
    .B(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4610_ (.B(_1424_),
    .A(_1391_),
    .X(_1425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4611_ (.Y(_1426_),
    .B(_1425_),
    .A_N(_1422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4612_ (.Y(_1427_),
    .A(_1422_),
    .B(_1425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4613_ (.B1(_1399_),
    .VDD(VPWR),
    .Y(_1428_),
    .VSS(VGND),
    .A1(_1397_),
    .A2(_1400_));
 sg13g2_nand2_1 _4614_ (.Y(_1429_),
    .A(net827),
    .B(net878),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4615_ (.A(net835),
    .B(net832),
    .C(net876),
    .D(net874),
    .X(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4616_ (.B(net831),
    .C(net876),
    .A(net836),
    .Y(_1431_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net874));
 sg13g2_a22oi_1 _4617_ (.Y(_1432_),
    .B1(net874),
    .B2(net836),
    .A2(net876),
    .A1(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4618_ (.A(_1429_),
    .B(_1430_),
    .C(_1432_),
    .X(_1433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4619_ (.B1(_1429_),
    .VDD(VPWR),
    .Y(_1434_),
    .VSS(VGND),
    .A1(_1430_),
    .A2(_1432_));
 sg13g2_and3_1 _4620_ (.X(_1435_),
    .A(_1428_),
    .B(_1433_),
    .C(_1434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4621_ (.B(_1433_),
    .C(_1434_),
    .A(_1428_),
    .Y(_1436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4622_ (.A2(_1434_),
    .A1(_1433_),
    .B1(_1428_),
    .X(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4623_ (.B(_1436_),
    .C(_1437_),
    .A(_1427_),
    .Y(_1438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4624_ (.A2(_1437_),
    .A1(_1436_),
    .B1(_1427_),
    .X(_1439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4625_ (.B(_1438_),
    .C(_1439_),
    .A(_1421_),
    .Y(_1440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4626_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1438_),
    .A2(_1439_),
    .Y(_1441_),
    .B1(_1421_));
 sg13g2_a21o_1 _4627_ (.A2(_1439_),
    .A1(_1438_),
    .B1(_1421_),
    .X(_1442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4628_ (.Y(_1443_),
    .A(_1440_),
    .B(_1442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4629_ (.Y(_1444_),
    .A(_1420_),
    .B(_1443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4630_ (.Y(_1445_),
    .B(_1416_),
    .A_N(_1444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4631_ (.B(_1444_),
    .A(_1416_),
    .X(_1446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4632_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1388_),
    .A2(_1414_),
    .Y(_1447_),
    .B1(_1413_));
 sg13g2_xor2_1 _4633_ (.B(_1447_),
    .A(_1446_),
    .X(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4634_ (.B1(_1440_),
    .VDD(VPWR),
    .Y(_1448_),
    .VSS(VGND),
    .A1(_1420_),
    .A2(_1441_));
 sg13g2_o21ai_1 _4635_ (.B1(_1426_),
    .VDD(VPWR),
    .Y(_1449_),
    .VSS(VGND),
    .A1(_1391_),
    .A2(_1424_));
 sg13g2_a22oi_1 _4636_ (.Y(_1450_),
    .B1(net820),
    .B2(\DP_3.matrix[0] ),
    .A2(net821),
    .A1(net885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4637_ (.Y(_1451_),
    .A(net885),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4638_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1452_),
    .B(_1451_),
    .A(_1418_));
 sg13g2_nor2b_1 _4639_ (.A(_1450_),
    .B_N(_1452_),
    .Y(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4640_ (.A(_1449_),
    .B(_1453_),
    .X(_1454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4641_ (.Y(_1455_),
    .A(_1449_),
    .B(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4642_ (.A2(_1437_),
    .A1(_1427_),
    .B1(_1435_),
    .X(_1456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4643_ (.Y(_1457_),
    .A(net883),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4644_ (.Y(_1458_),
    .A(net826),
    .B(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4645_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1459_),
    .B(_1458_),
    .A(_1423_));
 sg13g2_xnor2_1 _4646_ (.Y(_1460_),
    .A(_1423_),
    .B(_1458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4647_ (.Y(_1461_),
    .A(_1457_),
    .B(_1460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4648_ (.B1(_1431_),
    .VDD(VPWR),
    .Y(_1462_),
    .VSS(VGND),
    .A1(_1429_),
    .A2(_1432_));
 sg13g2_nand2_1 _4649_ (.Y(_1463_),
    .A(net827),
    .B(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4650_ (.A(net835),
    .B(net831),
    .C(net874),
    .D(net873),
    .X(_1464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4651_ (.B(net831),
    .C(net874),
    .A(net835),
    .Y(_1465_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net873));
 sg13g2_a22oi_1 _4652_ (.Y(_1466_),
    .B1(net873),
    .B2(net836),
    .A2(net874),
    .A1(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4653_ (.A(_1463_),
    .B(_1464_),
    .C(_1466_),
    .X(_1467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4654_ (.B1(_1463_),
    .VDD(VPWR),
    .Y(_1468_),
    .VSS(VGND),
    .A1(_1464_),
    .A2(_1466_));
 sg13g2_and3_1 _4655_ (.X(_1469_),
    .A(_1462_),
    .B(_1467_),
    .C(_1468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4656_ (.B(_1467_),
    .C(_1468_),
    .A(_1462_),
    .Y(_1470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4657_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1467_),
    .A2(_1468_),
    .Y(_1471_),
    .B1(_1462_));
 sg13g2_or3_1 _4658_ (.A(_1461_),
    .B(_1469_),
    .C(_1471_),
    .X(_1472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4659_ (.B1(_1461_),
    .VDD(VPWR),
    .Y(_1473_),
    .VSS(VGND),
    .A1(_1469_),
    .A2(_1471_));
 sg13g2_and3_1 _4660_ (.X(_1474_),
    .A(_1456_),
    .B(_1472_),
    .C(_1473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4661_ (.B(_1472_),
    .C(_1473_),
    .A(_1456_),
    .Y(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4662_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1472_),
    .A2(_1473_),
    .Y(_1476_),
    .B1(_1456_));
 sg13g2_or3_1 _4663_ (.A(_1455_),
    .B(_1474_),
    .C(_1476_),
    .X(_1477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4664_ (.B1(_1455_),
    .VDD(VPWR),
    .Y(_1478_),
    .VSS(VGND),
    .A1(_1474_),
    .A2(_1476_));
 sg13g2_nand3_1 _4665_ (.B(_1477_),
    .C(_1478_),
    .A(_1448_),
    .Y(_1479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1477_),
    .A2(_1478_),
    .Y(_1480_),
    .B1(_1448_));
 sg13g2_a21o_1 _4667_ (.A2(_1478_),
    .A1(_1477_),
    .B1(_1448_),
    .X(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4668_ (.Y(_1482_),
    .A(_1479_),
    .B(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4669_ (.B(_1482_),
    .A(_1419_),
    .X(_1483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4670_ (.B1(_1445_),
    .VDD(VPWR),
    .Y(_1484_),
    .VSS(VGND),
    .A1(_1446_),
    .A2(_1447_));
 sg13g2_nand2_1 _4671_ (.Y(_1485_),
    .A(_1483_),
    .B(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4672_ (.B(_1484_),
    .A(_1483_),
    .X(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4673_ (.B1(_1475_),
    .VDD(VPWR),
    .Y(_1486_),
    .VSS(VGND),
    .A1(_1455_),
    .A2(_1476_));
 sg13g2_o21ai_1 _4674_ (.B1(_1459_),
    .VDD(VPWR),
    .Y(_1487_),
    .VSS(VGND),
    .A1(_1457_),
    .A2(_1460_));
 sg13g2_nand2_1 _4675_ (.Y(_1488_),
    .A(\DP_3.matrix[0] ),
    .B(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4676_ (.Y(_1489_),
    .A(net883),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4677_ (.Y(_1490_),
    .A(net883),
    .B(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4678_ (.B(_1490_),
    .A(_1451_),
    .X(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4679_ (.Y(_1492_),
    .B(_1491_),
    .A_N(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4680_ (.Y(_1493_),
    .A(_1488_),
    .B(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4681_ (.Y(_1494_),
    .A(_1487_),
    .B(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4682_ (.Y(_1495_),
    .A(_1487_),
    .B(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4683_ (.Y(_1496_),
    .A(_1452_),
    .B(_1495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4684_ (.B1(_1470_),
    .VDD(VPWR),
    .Y(_1497_),
    .VSS(VGND),
    .A1(_1461_),
    .A2(_1471_));
 sg13g2_nand2_1 _4685_ (.Y(_1498_),
    .A(net881),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4686_ (.Y(_1499_),
    .A(net823),
    .B(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4687_ (.A(net825),
    .B(net879),
    .C(net823),
    .D(net877),
    .X(_1500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4688_ (.Y(_1501_),
    .B1(net877),
    .B2(net826),
    .A2(net823),
    .A1(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4689_ (.A(_1498_),
    .B(_1500_),
    .C(_1501_),
    .Y(_1502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4690_ (.B1(_1498_),
    .VDD(VPWR),
    .Y(_1503_),
    .VSS(VGND),
    .A1(_1500_),
    .A2(_1501_));
 sg13g2_nand2b_1 _4691_ (.Y(_1504_),
    .B(_1503_),
    .A_N(_1502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4692_ (.B1(_1465_),
    .VDD(VPWR),
    .Y(_1505_),
    .VSS(VGND),
    .A1(_1463_),
    .A2(_1466_));
 sg13g2_nand2_1 _4693_ (.Y(_1506_),
    .A(net828),
    .B(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4694_ (.A(net835),
    .B(net832),
    .C(net873),
    .D(net1001),
    .X(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4695_ (.B(net831),
    .C(net873),
    .A(net836),
    .Y(_1508_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1001));
 sg13g2_a22oi_1 _4696_ (.Y(_1509_),
    .B1(net1001),
    .B2(net835),
    .A2(net873),
    .A1(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4697_ (.A(_1506_),
    .B(_1507_),
    .C(_1509_),
    .X(_1510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4698_ (.B1(_1506_),
    .VDD(VPWR),
    .Y(_1511_),
    .VSS(VGND),
    .A1(_1507_),
    .A2(_1509_));
 sg13g2_and3_1 _4699_ (.X(_1512_),
    .A(_1505_),
    .B(_1510_),
    .C(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4700_ (.B(_1510_),
    .C(_1511_),
    .A(_1505_),
    .Y(_1513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1510_),
    .A2(_1511_),
    .Y(_1514_),
    .B1(_1505_));
 sg13g2_or3_1 _4702_ (.A(_1504_),
    .B(_1512_),
    .C(_1514_),
    .X(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4703_ (.B1(_1504_),
    .VDD(VPWR),
    .Y(_1516_),
    .VSS(VGND),
    .A1(_1512_),
    .A2(_1514_));
 sg13g2_and3_1 _4704_ (.X(_1517_),
    .A(_1497_),
    .B(_1515_),
    .C(_1516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4705_ (.B(_1515_),
    .C(_1516_),
    .A(_1497_),
    .Y(_1518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4706_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1515_),
    .A2(_1516_),
    .Y(_1519_),
    .B1(_1497_));
 sg13g2_or3_1 _4707_ (.A(_1496_),
    .B(_1517_),
    .C(_1519_),
    .X(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4708_ (.B1(_1496_),
    .VDD(VPWR),
    .Y(_1521_),
    .VSS(VGND),
    .A1(_1517_),
    .A2(_1519_));
 sg13g2_nand3_1 _4709_ (.B(_1520_),
    .C(_1521_),
    .A(_1486_),
    .Y(_1522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4710_ (.A2(_1521_),
    .A1(_1520_),
    .B1(_1486_),
    .X(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4711_ (.A2(_1523_),
    .A1(_1522_),
    .B1(_1454_),
    .X(_1524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4712_ (.B(_1522_),
    .C(_1523_),
    .A(_1454_),
    .Y(_1525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4713_ (.B1(_1479_),
    .VDD(VPWR),
    .Y(_1526_),
    .VSS(VGND),
    .A1(_1419_),
    .A2(_1480_));
 sg13g2_nand3_1 _4714_ (.B(_1525_),
    .C(_1526_),
    .A(_1524_),
    .Y(_1527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4715_ (.A2(_1525_),
    .A1(_1524_),
    .B1(_1526_),
    .X(_1528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4716_ (.A(_1527_),
    .B(_1528_),
    .X(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4717_ (.B(_1484_),
    .C(_1529_),
    .A(_1483_),
    .Y(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4718_ (.Y(_0147_),
    .A(_1485_),
    .B(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4719_ (.B1(_1494_),
    .VDD(VPWR),
    .Y(_1531_),
    .VSS(VGND),
    .A1(_1452_),
    .A2(_1495_));
 sg13g2_o21ai_1 _4720_ (.B1(_1518_),
    .VDD(VPWR),
    .Y(_1532_),
    .VSS(VGND),
    .A1(_1496_),
    .A2(_1519_));
 sg13g2_o21ai_1 _4721_ (.B1(_1492_),
    .VDD(VPWR),
    .Y(_1533_),
    .VSS(VGND),
    .A1(_1451_),
    .A2(_1490_));
 sg13g2_or2_1 _4722_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1534_),
    .B(_1502_),
    .A(_1500_));
 sg13g2_nand2_1 _4723_ (.Y(_1535_),
    .A(net885),
    .B(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4724_ (.Y(_1536_),
    .A(net881),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4725_ (.Y(_1537_),
    .A(net881),
    .B(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4726_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1538_),
    .B(_1536_),
    .A(_1490_));
 sg13g2_xnor2_1 _4727_ (.Y(_1539_),
    .A(_1489_),
    .B(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4728_ (.B(_1539_),
    .A(_1535_),
    .X(_1540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4729_ (.Y(_1541_),
    .A(_1534_),
    .B(_1540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4730_ (.A(_1541_),
    .B_N(_1533_),
    .Y(_1542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4731_ (.B(_1541_),
    .A(_1533_),
    .X(_1543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4732_ (.B1(_1513_),
    .VDD(VPWR),
    .Y(_1544_),
    .VSS(VGND),
    .A1(_1504_),
    .A2(_1514_));
 sg13g2_nand2_1 _4733_ (.Y(_1545_),
    .A(net879),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4734_ (.Y(_1546_),
    .A(net826),
    .B(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4735_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1547_),
    .B(_1546_),
    .A(_1499_));
 sg13g2_and2_1 _4736_ (.A(_1499_),
    .B(_1546_),
    .X(_1548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4737_ (.Y(_1549_),
    .A(_1499_),
    .B(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4738_ (.Y(_1550_),
    .A(_1545_),
    .B(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4739_ (.B1(_1508_),
    .VDD(VPWR),
    .Y(_1551_),
    .VSS(VGND),
    .A1(_1506_),
    .A2(_1509_));
 sg13g2_nand2_1 _4740_ (.Y(_1552_),
    .A(net828),
    .B(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4741_ (.A(net832),
    .B(net828),
    .C(net872),
    .D(net1002),
    .X(_1553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4742_ (.Y(_1554_),
    .B1(net1001),
    .B2(net831),
    .A2(net872),
    .A1(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4743_ (.A(_1553_),
    .B(_1554_),
    .Y(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4744_ (.Y(_1556_),
    .A(_1551_),
    .B(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4745_ (.Y(_1557_),
    .A(_1551_),
    .B(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4746_ (.B(_1557_),
    .A(_1550_),
    .X(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4747_ (.Y(_1559_),
    .A(_1544_),
    .B(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4748_ (.Y(_1560_),
    .A(_1544_),
    .B(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4749_ (.B(_1560_),
    .A(_1543_),
    .X(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4750_ (.Y(_1562_),
    .A(_1532_),
    .B(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4751_ (.Y(_1563_),
    .A(_1532_),
    .B(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4752_ (.Y(_1564_),
    .B(_1531_),
    .A_N(_1563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4753_ (.B(_1563_),
    .A(_1531_),
    .X(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4754_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1522_),
    .A2(_1525_),
    .Y(_1566_),
    .B1(_1565_));
 sg13g2_a21o_1 _4755_ (.A2(_1525_),
    .A1(_1522_),
    .B1(_1565_),
    .X(_1567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4756_ (.X(_1568_),
    .A(_1522_),
    .B(_1525_),
    .C(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4757_ (.A(_1566_),
    .B(_1568_),
    .Y(_1569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4758_ (.Y(_1570_),
    .A(_1527_),
    .B(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4759_ (.B(_1570_),
    .A(_1569_),
    .X(_0148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4760_ (.A2(_1540_),
    .A1(_1534_),
    .B1(_1542_),
    .X(_1571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4761_ (.B1(_1559_),
    .VDD(VPWR),
    .Y(_1572_),
    .VSS(VGND),
    .A1(_1543_),
    .A2(_1560_));
 sg13g2_o21ai_1 _4762_ (.B1(_1538_),
    .VDD(VPWR),
    .Y(_1573_),
    .VSS(VGND),
    .A1(_1535_),
    .A2(_1539_));
 sg13g2_o21ai_1 _4763_ (.B1(_1547_),
    .VDD(VPWR),
    .Y(_1574_),
    .VSS(VGND),
    .A1(_1545_),
    .A2(_1548_));
 sg13g2_nand2_1 _4764_ (.Y(_1575_),
    .A(net883),
    .B(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4765_ (.Y(_1576_),
    .A(net879),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4766_ (.Y(_1577_),
    .A(net879),
    .B(\DP_4.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4767_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1578_),
    .B(_1576_),
    .A(_1537_));
 sg13g2_xnor2_1 _4768_ (.Y(_1579_),
    .A(_1536_),
    .B(_1577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4769_ (.B(_1579_),
    .A(_1575_),
    .X(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4770_ (.Y(_1581_),
    .A(_1574_),
    .B(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4771_ (.A(_1581_),
    .B_N(_1573_),
    .Y(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4772_ (.B(_1581_),
    .A(_1573_),
    .X(_1583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4773_ (.B1(_1556_),
    .VDD(VPWR),
    .Y(_1584_),
    .VSS(VGND),
    .A1(_1550_),
    .A2(_1557_));
 sg13g2_a21oi_1 _4774_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net831),
    .A2(net872),
    .Y(_1585_),
    .B1(_1552_));
 sg13g2_nand2_1 _4775_ (.Y(_1586_),
    .A(net877),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4776_ (.Y(_1587_),
    .A(net823),
    .B(net872),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4777_ (.A(net825),
    .B(net823),
    .C(net875),
    .D(\DP_3.matrix[7] ),
    .X(_1588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4778_ (.Y(_1589_),
    .B1(net872),
    .B2(net826),
    .A2(net875),
    .A1(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4779_ (.A(_1586_),
    .B(_1588_),
    .C(_1589_),
    .Y(_1590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4780_ (.B1(_1586_),
    .VDD(VPWR),
    .Y(_1591_),
    .VSS(VGND),
    .A1(_1588_),
    .A2(_1589_));
 sg13g2_nor2b_1 _4781_ (.A(_1590_),
    .B_N(_1591_),
    .Y(_1592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4782_ (.Y(_1593_),
    .A(_1585_),
    .B(_1592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4783_ (.Y(_1594_),
    .B(_1584_),
    .A_N(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4784_ (.B(_1593_),
    .A(_1584_),
    .X(_1595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4785_ (.B(_1595_),
    .A(_1583_),
    .X(_1596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4786_ (.Y(_1597_),
    .A(_1572_),
    .B(_1596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4787_ (.B(_1596_),
    .A(_1572_),
    .X(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4788_ (.Y(_1599_),
    .A(_1571_),
    .B(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4789_ (.Y(_1600_),
    .A(_1571_),
    .B(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1562_),
    .A2(_1564_),
    .Y(_1601_),
    .B1(_1600_));
 sg13g2_nand3_1 _4791_ (.B(_1564_),
    .C(_1600_),
    .A(_1562_),
    .Y(_1602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4792_ (.A(_1601_),
    .B_N(_1602_),
    .Y(_1603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4793_ (.B(_1484_),
    .C(_1529_),
    .A(_1483_),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1569_));
 sg13g2_a21oi_1 _4794_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1527_),
    .A2(_1567_),
    .Y(_1605_),
    .B1(_1568_));
 sg13g2_nand2b_1 _4795_ (.Y(_1606_),
    .B(_1604_),
    .A_N(_1605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4796_ (.B(_1606_),
    .A(_1603_),
    .X(_0139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4797_ (.A2(_1580_),
    .A1(_1574_),
    .B1(_1582_),
    .X(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4798_ (.B1(_1594_),
    .VDD(VPWR),
    .Y(_1608_),
    .VSS(VGND),
    .A1(_1583_),
    .A2(_1595_));
 sg13g2_a21o_2 _4799_ (.A2(_1592_),
    .A1(_1585_),
    .B1(_1553_),
    .X(_1609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4800_ (.Y(_1610_),
    .A(\DP_4.matrix[5] ),
    .B(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4801_ (.Y(_1611_),
    .A(net826),
    .B(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4802_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1612_),
    .B(_1611_),
    .A(_1587_));
 sg13g2_xnor2_1 _4803_ (.Y(_1613_),
    .A(_1587_),
    .B(_1611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4804_ (.B(_1613_),
    .A(_1610_),
    .X(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4805_ (.Y(_1615_),
    .A(_1609_),
    .B(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4806_ (.B1(_1578_),
    .VDD(VPWR),
    .Y(_1616_),
    .VSS(VGND),
    .A1(_1575_),
    .A2(_1579_));
 sg13g2_or2_1 _4807_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1617_),
    .B(_1590_),
    .A(_1588_));
 sg13g2_nand2_1 _4808_ (.Y(_1618_),
    .A(net881),
    .B(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4809_ (.Y(_1619_),
    .A(net877),
    .B(\DP_4.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4810_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1620_),
    .B(_1619_),
    .A(_1576_));
 sg13g2_xnor2_1 _4811_ (.Y(_1621_),
    .A(_1576_),
    .B(_1619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4812_ (.B(_1621_),
    .A(_1618_),
    .X(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4813_ (.Y(_1623_),
    .A(_1617_),
    .B(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4814_ (.A(_1623_),
    .B_N(_1616_),
    .Y(_1624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4815_ (.B(_1623_),
    .A(_1616_),
    .X(_1625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4816_ (.A(_1615_),
    .B(_1625_),
    .Y(_1626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4817_ (.B(_1625_),
    .A(_1615_),
    .X(_1627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4818_ (.Y(_1628_),
    .A(_1608_),
    .B(_1627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4819_ (.A(_1628_),
    .B_N(_1607_),
    .Y(_1629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4820_ (.B(_1628_),
    .A(_1607_),
    .X(_1630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4821_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1597_),
    .A2(_1599_),
    .Y(_1631_),
    .B1(_1630_));
 sg13g2_nand3_1 _4822_ (.B(_1599_),
    .C(_1630_),
    .A(_1597_),
    .Y(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4823_ (.A(_1631_),
    .B_N(_1632_),
    .Y(_1633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4824_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1603_),
    .A2(_1606_),
    .Y(_1634_),
    .B1(_1601_));
 sg13g2_xnor2_1 _4825_ (.Y(_0140_),
    .A(_1633_),
    .B(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4826_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1617_),
    .A2(_1622_),
    .Y(_1635_),
    .B1(_1624_));
 sg13g2_a22oi_1 _4827_ (.Y(_1636_),
    .B1(net1002),
    .B2(net824),
    .A2(net872),
    .A1(\DP_4.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4828_ (.Y(_1637_),
    .A(\DP_4.matrix[5] ),
    .B(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4829_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1638_),
    .B(_1637_),
    .A(_1587_));
 sg13g2_nand2b_1 _4830_ (.Y(_1639_),
    .B(_1638_),
    .A_N(_1636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4831_ (.B1(_1620_),
    .VDD(VPWR),
    .Y(_1640_),
    .VSS(VGND),
    .A1(_1618_),
    .A2(_1621_));
 sg13g2_o21ai_1 _4832_ (.B1(_1612_),
    .VDD(VPWR),
    .Y(_1641_),
    .VSS(VGND),
    .A1(_1610_),
    .A2(_1613_));
 sg13g2_nand2_1 _4833_ (.Y(_1642_),
    .A(\DP_3.matrix[4] ),
    .B(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4834_ (.Y(_1643_),
    .A(net875),
    .B(\DP_4.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4835_ (.A(_1619_),
    .B(_1643_),
    .Y(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4836_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1645_),
    .B(_1643_),
    .A(_1619_));
 sg13g2_a22oi_1 _4837_ (.Y(_1646_),
    .B1(\DP_4.matrix[7] ),
    .B2(net877),
    .A2(net821),
    .A1(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4838_ (.A(_1644_),
    .B(_1646_),
    .Y(_1647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4839_ (.Y(_1648_),
    .A(_1642_),
    .B(_1647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4840_ (.Y(_1649_),
    .A(_1641_),
    .B(_1648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4841_ (.A(_1649_),
    .B_N(_1640_),
    .Y(_1650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4842_ (.B(_1649_),
    .A(_1640_),
    .X(_1651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4843_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1652_),
    .B(_1651_),
    .A(_1639_));
 sg13g2_xor2_1 _4844_ (.B(_1651_),
    .A(_1639_),
    .X(_1653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4845_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1609_),
    .A2(_1614_),
    .Y(_1654_),
    .B1(_1626_));
 sg13g2_nand2b_1 _4846_ (.Y(_1655_),
    .B(_1653_),
    .A_N(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4847_ (.A(_1653_),
    .B_N(_1654_),
    .Y(_1656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4848_ (.B(_1654_),
    .A(_1653_),
    .X(_1657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4849_ (.Y(_1658_),
    .A(_1635_),
    .B(_1657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1608_),
    .A2(_1627_),
    .Y(_1659_),
    .B1(_1629_));
 sg13g2_or2_1 _4851_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1660_),
    .B(_1659_),
    .A(_1658_));
 sg13g2_xor2_1 _4852_ (.B(_1659_),
    .A(_1658_),
    .X(_1661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4853_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1601_),
    .A2(_1632_),
    .Y(_1662_),
    .B1(_1631_));
 sg13g2_nor2b_1 _4854_ (.A(_1605_),
    .B_N(_1662_),
    .Y(_1663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4855_ (.B1(_1632_),
    .VDD(VPWR),
    .Y(_1664_),
    .VSS(VGND),
    .A1(_1602_),
    .A2(_1631_));
 sg13g2_a21oi_2 _4856_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1664_),
    .Y(_1665_),
    .A2(_1663_),
    .A1(_1604_));
 sg13g2_nand2_1 _4857_ (.Y(_1666_),
    .A(_1661_),
    .B(_1665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4858_ (.B(_1665_),
    .A(_1661_),
    .X(_0141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4859_ (.B1(_1655_),
    .VDD(VPWR),
    .Y(_1667_),
    .VSS(VGND),
    .A1(_1635_),
    .A2(_1656_));
 sg13g2_a21o_1 _4860_ (.A2(_1648_),
    .A1(_1641_),
    .B1(_1650_),
    .X(_1668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4861_ (.B1(_1645_),
    .VDD(VPWR),
    .Y(_1669_),
    .VSS(VGND),
    .A1(_1642_),
    .A2(_1646_));
 sg13g2_nand2_1 _4862_ (.Y(_1670_),
    .A(net877),
    .B(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4863_ (.Y(_1671_),
    .A(net872),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4864_ (.Y(_1672_),
    .A(net821),
    .B(\DP_3.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4865_ (.B(_1672_),
    .A(_1643_),
    .X(_1673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4866_ (.Y(_1674_),
    .B(_1673_),
    .A_N(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4867_ (.Y(_1675_),
    .A(_1670_),
    .B(_1673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4868_ (.A(_1638_),
    .B_N(_1675_),
    .Y(_1676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4869_ (.Y(_1677_),
    .A(_1638_),
    .B(_1675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4870_ (.Y(_1678_),
    .A(_1669_),
    .B(_1677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4871_ (.A(_1637_),
    .B(_1678_),
    .Y(_1679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4872_ (.B(_1678_),
    .A(_1637_),
    .X(_1680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4873_ (.Y(_1681_),
    .B(_1680_),
    .A_N(_1652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4874_ (.Y(_1682_),
    .A(_1652_),
    .B(_1680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4875_ (.Y(_1683_),
    .A(_1668_),
    .B(_1682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4876_ (.B(_1682_),
    .A(_1668_),
    .X(_1684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4877_ (.A(_1667_),
    .B(_1684_),
    .Y(_1685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4878_ (.Y(_1686_),
    .A(_1667_),
    .B(_1684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4879_ (.A(_1685_),
    .B_N(_1686_),
    .Y(_1687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4880_ (.Y(_1688_),
    .A(_1660_),
    .B(_1666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4881_ (.B(_1688_),
    .A(_1687_),
    .X(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4882_ (.A(_1661_),
    .B(_1687_),
    .X(_1689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4883_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1660_),
    .A2(_1686_),
    .Y(_1690_),
    .B1(_1685_));
 sg13g2_a21o_1 _4884_ (.A2(_1689_),
    .A1(_1665_),
    .B1(_1690_),
    .X(_1691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4885_ (.A(_1681_),
    .B(_1683_),
    .X(_1692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4886_ (.A2(_1677_),
    .A1(_1669_),
    .B1(_1676_),
    .X(_1693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4887_ (.Y(_1694_),
    .A(net875),
    .B(\DP_4.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4888_ (.Y(_1695_),
    .A(\DP_4.matrix[7] ),
    .B(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4889_ (.Y(_1696_),
    .A(\DP_4.matrix[6] ),
    .B(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4890_ (.B(_1696_),
    .A(_1671_),
    .X(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4891_ (.Y(_1698_),
    .B(_1697_),
    .A_N(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4892_ (.Y(_1699_),
    .A(_1694_),
    .B(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4893_ (.B1(_1674_),
    .VDD(VPWR),
    .Y(_1700_),
    .VSS(VGND),
    .A1(_1643_),
    .A2(_1672_));
 sg13g2_nand2_1 _4894_ (.Y(_1701_),
    .A(_1699_),
    .B(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4895_ (.B(_1700_),
    .A(_1699_),
    .X(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4896_ (.Y(_1703_),
    .A(_1679_),
    .B(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4897_ (.A(_1703_),
    .B_N(_1693_),
    .Y(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4898_ (.B(_1703_),
    .A(_1693_),
    .X(_1705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4899_ (.A(_1692_),
    .B(_1705_),
    .Y(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4900_ (.B(_1705_),
    .A(_1692_),
    .X(_1707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4901_ (.B(_1707_),
    .A(_1691_),
    .X(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4902_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1691_),
    .A2(_1707_),
    .Y(_1708_),
    .B1(_1706_));
 sg13g2_a21oi_1 _4903_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1679_),
    .A2(_1702_),
    .Y(_1709_),
    .B1(_1704_));
 sg13g2_o21ai_1 _4904_ (.B1(_1698_),
    .VDD(VPWR),
    .Y(_1710_),
    .VSS(VGND),
    .A1(_1671_),
    .A2(_1696_));
 sg13g2_nand2_1 _4905_ (.Y(_1711_),
    .A(net872),
    .B(\DP_4.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4906_ (.Y(_1712_),
    .A(_1695_),
    .B(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4907_ (.Y(_1713_),
    .A(_1710_),
    .B(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4908_ (.Y(_1714_),
    .A(_1701_),
    .B(_1713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4909_ (.Y(_1715_),
    .A(_1709_),
    .B(_1714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4910_ (.Y(_0144_),
    .A(_1708_),
    .B(_1715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4911_ (.A(net279),
    .B(net800),
    .X(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4912_ (.X(_1716_),
    .A(net853),
    .B(net796),
    .C(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4913_ (.Y(_1717_),
    .B1(net796),
    .B2(net279),
    .A2(net853),
    .A1(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4914_ (.A(_1716_),
    .B(net289),
    .Y(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4915_ (.A(net854),
    .B(net792),
    .X(_1718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4916_ (.A(net799),
    .B(net853),
    .C(net796),
    .D(net851),
    .X(_1719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4917_ (.Y(_1720_),
    .B1(net851),
    .B2(net799),
    .A2(net796),
    .A1(net853),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4918_ (.A(_1719_),
    .B(_1720_),
    .Y(_1721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4919_ (.B(_1721_),
    .A(_1718_),
    .X(_1722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4920_ (.Y(_1723_),
    .A(_1716_),
    .B(_1722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4921_ (.B(_1722_),
    .A(_1716_),
    .X(_0091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4922_ (.Y(_1724_),
    .A(net854),
    .B(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4923_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1718_),
    .A2(_1721_),
    .Y(_1725_),
    .B1(_1719_));
 sg13g2_nand2_1 _4924_ (.Y(_1726_),
    .A(net852),
    .B(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4925_ (.A(net799),
    .B(net795),
    .C(net851),
    .D(net848),
    .X(_1727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4926_ (.B(\DP_4.matrix[73] ),
    .C(net851),
    .A(net799),
    .Y(_1728_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net848));
 sg13g2_a22oi_1 _4927_ (.Y(_1729_),
    .B1(net849),
    .B2(net799),
    .A2(net850),
    .A1(\DP_4.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4928_ (.A(_1726_),
    .B(_1727_),
    .C(_1729_),
    .Y(_1730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4929_ (.B1(_1726_),
    .VDD(VPWR),
    .Y(_1731_),
    .VSS(VGND),
    .A1(_1727_),
    .A2(_1729_));
 sg13g2_nor2b_1 _4930_ (.A(_1730_),
    .B_N(_1731_),
    .Y(_1732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4931_ (.Y(_1733_),
    .B(_1732_),
    .A_N(_1725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4932_ (.Y(_1734_),
    .A(_1725_),
    .B(_1732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4933_ (.Y(_1735_),
    .B(_1734_),
    .A_N(_1724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4934_ (.Y(_1736_),
    .A(_1724_),
    .B(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4935_ (.A(_1723_),
    .B_N(_1736_),
    .Y(_1737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4936_ (.Y(_0092_),
    .A(_1723_),
    .B(_1736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4937_ (.Y(_1738_),
    .B1(net787),
    .B2(net854),
    .A2(net789),
    .A1(net852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4938_ (.Y(_1739_),
    .A(net852),
    .B(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4939_ (.A(_1724_),
    .B(_1739_),
    .Y(_1740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4940_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1741_),
    .B(_1740_),
    .A(_1738_));
 sg13g2_o21ai_1 _4941_ (.B1(_1728_),
    .VDD(VPWR),
    .Y(_1742_),
    .VSS(VGND),
    .A1(_1726_),
    .A2(_1729_));
 sg13g2_nand2_1 _4942_ (.Y(_1743_),
    .A(net850),
    .B(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4943_ (.A(net799),
    .B(net795),
    .C(net849),
    .D(net847),
    .X(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4944_ (.B(net795),
    .C(net849),
    .A(net799),
    .Y(_1745_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net847));
 sg13g2_a22oi_1 _4945_ (.Y(_1746_),
    .B1(net847),
    .B2(net799),
    .A2(net849),
    .A1(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4946_ (.A(_1743_),
    .B(_1744_),
    .C(_1746_),
    .X(_1747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4947_ (.B1(_1743_),
    .VDD(VPWR),
    .Y(_1748_),
    .VSS(VGND),
    .A1(_1744_),
    .A2(_1746_));
 sg13g2_nand3_1 _4948_ (.B(_1747_),
    .C(_1748_),
    .A(_1742_),
    .Y(_1749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4949_ (.A2(_1748_),
    .A1(_1747_),
    .B1(_1742_),
    .X(_1750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4950_ (.Y(_1751_),
    .A(_1749_),
    .B(_1750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4951_ (.B(_1751_),
    .A(_1741_),
    .X(_1752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4952_ (.Y(_1753_),
    .A(_1733_),
    .B(_1735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4953_ (.Y(_1754_),
    .A(_1752_),
    .B(_1753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4954_ (.B(_1753_),
    .A(_1752_),
    .X(_1755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4955_ (.A(_1737_),
    .B(_1755_),
    .X(_1756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4956_ (.B(_1755_),
    .A(_1737_),
    .X(_0093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4957_ (.B1(_1749_),
    .VDD(VPWR),
    .Y(_1757_),
    .VSS(VGND),
    .A1(_1741_),
    .A2(_1751_));
 sg13g2_nand2_1 _4958_ (.Y(_1758_),
    .A(net854),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4959_ (.Y(_1759_),
    .A(net850),
    .B(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4960_ (.Y(_1760_),
    .A(net850),
    .B(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4961_ (.B(_1760_),
    .A(_1739_),
    .X(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4962_ (.Y(_1762_),
    .B(_1761_),
    .A_N(_1758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4963_ (.B(_1761_),
    .A(_1758_),
    .X(_1763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4964_ (.B1(_1745_),
    .VDD(VPWR),
    .Y(_1764_),
    .VSS(VGND),
    .A1(_1743_),
    .A2(_1746_));
 sg13g2_nand2_1 _4965_ (.Y(_1765_),
    .A(net791),
    .B(net849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4966_ (.A(net798),
    .B(net795),
    .C(net846),
    .D(net845),
    .X(_1766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4967_ (.B(net795),
    .C(net846),
    .A(net798),
    .Y(_1767_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net844));
 sg13g2_a22oi_1 _4968_ (.Y(_1768_),
    .B1(net845),
    .B2(net798),
    .A2(net847),
    .A1(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4969_ (.A(_1765_),
    .B(_1766_),
    .C(_1768_),
    .X(_1769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4970_ (.B1(_1765_),
    .VDD(VPWR),
    .Y(_1770_),
    .VSS(VGND),
    .A1(_1766_),
    .A2(_1768_));
 sg13g2_and3_1 _4971_ (.X(_1771_),
    .A(_1764_),
    .B(_1769_),
    .C(_1770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4972_ (.B(_1769_),
    .C(_1770_),
    .A(_1764_),
    .Y(_1772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4973_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1769_),
    .A2(_1770_),
    .Y(_1773_),
    .B1(_1764_));
 sg13g2_or3_1 _4974_ (.A(_1763_),
    .B(_1771_),
    .C(_1773_),
    .X(_1774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4975_ (.B1(_1763_),
    .VDD(VPWR),
    .Y(_1775_),
    .VSS(VGND),
    .A1(_1771_),
    .A2(_1773_));
 sg13g2_nand3_1 _4976_ (.B(_1774_),
    .C(_1775_),
    .A(_1757_),
    .Y(_1776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4977_ (.A2(_1775_),
    .A1(_1774_),
    .B1(_1757_),
    .X(_1777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1776_),
    .A2(_1777_),
    .Y(_1778_),
    .B1(_1740_));
 sg13g2_and3_1 _4979_ (.X(_1779_),
    .A(_1740_),
    .B(_1776_),
    .C(_1777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4980_ (.B(_1776_),
    .C(_1777_),
    .A(_1740_),
    .Y(_1780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4981_ (.A(_1754_),
    .B(_1778_),
    .C(_1779_),
    .Y(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4982_ (.B1(_1754_),
    .VDD(VPWR),
    .Y(_1782_),
    .VSS(VGND),
    .A1(_1778_),
    .A2(_1779_));
 sg13g2_nand2b_1 _4983_ (.Y(_1783_),
    .B(_1782_),
    .A_N(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4984_ (.Y(_0149_),
    .A(_1756_),
    .B(_1783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4985_ (.Y(_1784_),
    .A(_1776_),
    .B(_1780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4986_ (.B1(_1762_),
    .VDD(VPWR),
    .Y(_1785_),
    .VSS(VGND),
    .A1(_1739_),
    .A2(_1760_));
 sg13g2_nand2_1 _4987_ (.Y(_1786_),
    .A(net854),
    .B(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4988_ (.Y(_1787_),
    .B(_1785_),
    .A_N(_1786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4989_ (.B(_1786_),
    .A(_1785_),
    .X(_1788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4990_ (.B1(_1772_),
    .VDD(VPWR),
    .Y(_1789_),
    .VSS(VGND),
    .A1(_1763_),
    .A2(_1773_));
 sg13g2_nand2_1 _4991_ (.Y(_1790_),
    .A(net852),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4992_ (.Y(_1791_),
    .A(net848),
    .B(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4993_ (.Y(_1792_),
    .A(net848),
    .B(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4994_ (.B(_1792_),
    .A(_1759_),
    .X(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4995_ (.Y(_1794_),
    .B(_1793_),
    .A_N(_1790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4996_ (.Y(_1795_),
    .A(_1790_),
    .B(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4997_ (.B1(_1767_),
    .VDD(VPWR),
    .Y(_1796_),
    .VSS(VGND),
    .A1(_1765_),
    .A2(_1768_));
 sg13g2_nand2_1 _4998_ (.Y(_1797_),
    .A(net791),
    .B(net847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4999_ (.A(net797),
    .B(net793),
    .C(net844),
    .D(net841),
    .X(_1798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5000_ (.B(net793),
    .C(net845),
    .A(net797),
    .Y(_1799_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net842));
 sg13g2_a22oi_1 _5001_ (.Y(_1800_),
    .B1(net841),
    .B2(net797),
    .A2(net845),
    .A1(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5002_ (.A(_1797_),
    .B(_1798_),
    .C(_1800_),
    .X(_1801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5003_ (.B1(_1797_),
    .VDD(VPWR),
    .Y(_1802_),
    .VSS(VGND),
    .A1(_1798_),
    .A2(_1800_));
 sg13g2_and3_1 _5004_ (.X(_1803_),
    .A(_1796_),
    .B(_1801_),
    .C(_1802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5005_ (.B(_1801_),
    .C(_1802_),
    .A(_1796_),
    .Y(_1804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5006_ (.A2(_1802_),
    .A1(_1801_),
    .B1(_1796_),
    .X(_1805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5007_ (.B(_1804_),
    .C(_1805_),
    .A(_1795_),
    .Y(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5008_ (.A2(_1805_),
    .A1(_1804_),
    .B1(_1795_),
    .X(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5009_ (.B(_1806_),
    .C(_1807_),
    .A(_1789_),
    .Y(_1808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5010_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1806_),
    .A2(_1807_),
    .Y(_1809_),
    .B1(_1789_));
 sg13g2_a21o_1 _5011_ (.A2(_1807_),
    .A1(_1806_),
    .B1(_1789_),
    .X(_1810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5012_ (.Y(_1811_),
    .A(_1808_),
    .B(_1810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5013_ (.Y(_1812_),
    .A(_1788_),
    .B(_1811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5014_ (.Y(_1813_),
    .B(_1784_),
    .A_N(_1812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5015_ (.B(_1812_),
    .A(_1784_),
    .X(_1814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5016_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1756_),
    .A2(_1782_),
    .Y(_1815_),
    .B1(_1781_));
 sg13g2_xor2_1 _5017_ (.B(_1815_),
    .A(_1814_),
    .X(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5018_ (.B1(_1808_),
    .VDD(VPWR),
    .Y(_1816_),
    .VSS(VGND),
    .A1(_1788_),
    .A2(_1809_));
 sg13g2_o21ai_1 _5019_ (.B1(_1794_),
    .VDD(VPWR),
    .Y(_1817_),
    .VSS(VGND),
    .A1(_1759_),
    .A2(_1792_));
 sg13g2_a22oi_1 _5020_ (.Y(_1818_),
    .B1(net781),
    .B2(net854),
    .A2(net783),
    .A1(net852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5021_ (.Y(_1819_),
    .A(net852),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5022_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1820_),
    .B(_1819_),
    .A(_1786_));
 sg13g2_nor2b_1 _5023_ (.A(_1818_),
    .B_N(_1820_),
    .Y(_1821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5024_ (.A(_1817_),
    .B(_1821_),
    .X(_1822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5025_ (.Y(_1823_),
    .A(_1817_),
    .B(_1821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5026_ (.A2(_1805_),
    .A1(_1795_),
    .B1(_1803_),
    .X(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5027_ (.Y(_1825_),
    .A(net850),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5028_ (.Y(_1826_),
    .A(net846),
    .B(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5029_ (.Y(_1827_),
    .A(net789),
    .B(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5030_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1828_),
    .B(_1826_),
    .A(_1792_));
 sg13g2_xnor2_1 _5031_ (.Y(_1829_),
    .A(_1791_),
    .B(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5032_ (.Y(_1830_),
    .A(_1825_),
    .B(_1829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5033_ (.B1(_1799_),
    .VDD(VPWR),
    .Y(_1831_),
    .VSS(VGND),
    .A1(_1797_),
    .A2(_1800_));
 sg13g2_nand2_1 _5034_ (.Y(_1832_),
    .A(net791),
    .B(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5035_ (.A(net797),
    .B(net793),
    .C(net842),
    .D(net839),
    .X(_1833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5036_ (.B(net793),
    .C(net842),
    .A(net797),
    .Y(_1834_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net839));
 sg13g2_a22oi_1 _5037_ (.Y(_1835_),
    .B1(net839),
    .B2(net797),
    .A2(net842),
    .A1(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5038_ (.A(_1832_),
    .B(_1833_),
    .C(_1835_),
    .X(_1836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5039_ (.B1(_1832_),
    .VDD(VPWR),
    .Y(_1837_),
    .VSS(VGND),
    .A1(_1833_),
    .A2(_1835_));
 sg13g2_and3_1 _5040_ (.X(_1838_),
    .A(_1831_),
    .B(_1836_),
    .C(_1837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5041_ (.B(_1836_),
    .C(_1837_),
    .A(_1831_),
    .Y(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5042_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1836_),
    .A2(_1837_),
    .Y(_1840_),
    .B1(_1831_));
 sg13g2_or3_1 _5043_ (.A(_1830_),
    .B(_1838_),
    .C(_1840_),
    .X(_1841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5044_ (.B1(_1830_),
    .VDD(VPWR),
    .Y(_1842_),
    .VSS(VGND),
    .A1(_1838_),
    .A2(_1840_));
 sg13g2_and3_1 _5045_ (.X(_1843_),
    .A(_1824_),
    .B(_1841_),
    .C(_1842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5046_ (.B(_1841_),
    .C(_1842_),
    .A(_1824_),
    .Y(_1844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5047_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1841_),
    .A2(_1842_),
    .Y(_1845_),
    .B1(_1824_));
 sg13g2_or3_1 _5048_ (.A(_1823_),
    .B(_1843_),
    .C(_1845_),
    .X(_1846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5049_ (.B1(_1823_),
    .VDD(VPWR),
    .Y(_1847_),
    .VSS(VGND),
    .A1(_1843_),
    .A2(_1845_));
 sg13g2_nand3_1 _5050_ (.B(_1846_),
    .C(_1847_),
    .A(_1816_),
    .Y(_1848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5051_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1846_),
    .A2(_1847_),
    .Y(_1849_),
    .B1(_1816_));
 sg13g2_a21o_1 _5052_ (.A2(_1847_),
    .A1(_1846_),
    .B1(_1816_),
    .X(_1850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5053_ (.Y(_1851_),
    .A(_1848_),
    .B(_1850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5054_ (.B(_1851_),
    .A(_1787_),
    .X(_1852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5055_ (.B1(_1813_),
    .VDD(VPWR),
    .Y(_1853_),
    .VSS(VGND),
    .A1(_1814_),
    .A2(_1815_));
 sg13g2_nand2_1 _5056_ (.Y(_1854_),
    .A(_1852_),
    .B(_1853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5057_ (.B(_1853_),
    .A(_1852_),
    .X(_0157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5058_ (.B1(_1844_),
    .VDD(VPWR),
    .Y(_1855_),
    .VSS(VGND),
    .A1(_1823_),
    .A2(_1845_));
 sg13g2_o21ai_1 _5059_ (.B1(_1828_),
    .VDD(VPWR),
    .Y(_1856_),
    .VSS(VGND),
    .A1(_1825_),
    .A2(_1829_));
 sg13g2_nand2_1 _5060_ (.Y(_1857_),
    .A(net854),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5061_ (.Y(_1858_),
    .A(net850),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5062_ (.Y(_1859_),
    .A(net850),
    .B(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5063_ (.B(_1859_),
    .A(_1819_),
    .X(_1860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5064_ (.Y(_1861_),
    .B(_1860_),
    .A_N(_1857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5065_ (.Y(_1862_),
    .A(_1857_),
    .B(_1860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5066_ (.Y(_1863_),
    .A(_1856_),
    .B(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5067_ (.Y(_1864_),
    .A(_1856_),
    .B(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5068_ (.Y(_1865_),
    .A(_1820_),
    .B(_1864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5069_ (.B1(_1839_),
    .VDD(VPWR),
    .Y(_1866_),
    .VSS(VGND),
    .A1(_1830_),
    .A2(_1840_));
 sg13g2_nand2_1 _5070_ (.Y(_1867_),
    .A(net848),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5071_ (.Y(_1868_),
    .A(net787),
    .B(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5072_ (.Y(_1869_),
    .A(net789),
    .B(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5073_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1870_),
    .B(_1868_),
    .A(_1827_));
 sg13g2_and2_1 _5074_ (.A(_1826_),
    .B(_1869_),
    .X(_1871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5075_ (.Y(_1872_),
    .A(_1826_),
    .B(_1869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5076_ (.Y(_1873_),
    .A(_1867_),
    .B(_1872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5077_ (.B1(_1834_),
    .VDD(VPWR),
    .Y(_1874_),
    .VSS(VGND),
    .A1(_1832_),
    .A2(_1835_));
 sg13g2_nand2_1 _5078_ (.Y(_1875_),
    .A(net791),
    .B(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5079_ (.A(net797),
    .B(net794),
    .C(net839),
    .D(net997),
    .X(_1876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5080_ (.B(net793),
    .C(net839),
    .A(net798),
    .Y(_1877_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net998));
 sg13g2_a22oi_1 _5081_ (.Y(_1878_),
    .B1(net998),
    .B2(net797),
    .A2(net839),
    .A1(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5082_ (.A(_1875_),
    .B(_1876_),
    .C(_1878_),
    .X(_1879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5083_ (.B1(_1875_),
    .VDD(VPWR),
    .Y(_1880_),
    .VSS(VGND),
    .A1(_1876_),
    .A2(_1878_));
 sg13g2_and3_1 _5084_ (.X(_1881_),
    .A(_1874_),
    .B(_1879_),
    .C(_1880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5085_ (.B(_1879_),
    .C(_1880_),
    .A(_1874_),
    .Y(_1882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5086_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1879_),
    .A2(_1880_),
    .Y(_1883_),
    .B1(_1874_));
 sg13g2_or3_1 _5087_ (.A(_1873_),
    .B(_1881_),
    .C(_1883_),
    .X(_1884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5088_ (.B1(_1873_),
    .VDD(VPWR),
    .Y(_1885_),
    .VSS(VGND),
    .A1(_1881_),
    .A2(_1883_));
 sg13g2_and3_1 _5089_ (.X(_1886_),
    .A(_1866_),
    .B(_1884_),
    .C(_1885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5090_ (.B(_1884_),
    .C(_1885_),
    .A(_1866_),
    .Y(_1887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5091_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1884_),
    .A2(_1885_),
    .Y(_1888_),
    .B1(_1866_));
 sg13g2_or3_1 _5092_ (.A(_1865_),
    .B(_1886_),
    .C(_1888_),
    .X(_1889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5093_ (.B1(_1865_),
    .VDD(VPWR),
    .Y(_1890_),
    .VSS(VGND),
    .A1(_1886_),
    .A2(_1888_));
 sg13g2_nand3_1 _5094_ (.B(_1889_),
    .C(_1890_),
    .A(_1855_),
    .Y(_1891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5095_ (.A2(_1890_),
    .A1(_1889_),
    .B1(_1855_),
    .X(_1892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5096_ (.A2(_1892_),
    .A1(_1891_),
    .B1(_1822_),
    .X(_1893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5097_ (.B(_1891_),
    .C(_1892_),
    .A(_1822_),
    .Y(_1894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5098_ (.B1(_1848_),
    .VDD(VPWR),
    .Y(_1895_),
    .VSS(VGND),
    .A1(_1787_),
    .A2(_1849_));
 sg13g2_nand3_1 _5099_ (.B(_1894_),
    .C(_1895_),
    .A(_1893_),
    .Y(_1896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5100_ (.A2(_1894_),
    .A1(_1893_),
    .B1(_1895_),
    .X(_1897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5101_ (.A(_1896_),
    .B(_1897_),
    .X(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5102_ (.B(_1853_),
    .C(_1898_),
    .A(_1852_),
    .Y(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5103_ (.Y(_0158_),
    .A(_1854_),
    .B(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5104_ (.B1(_1863_),
    .VDD(VPWR),
    .Y(_1900_),
    .VSS(VGND),
    .A1(_1820_),
    .A2(_1864_));
 sg13g2_o21ai_1 _5105_ (.B1(_1887_),
    .VDD(VPWR),
    .Y(_1901_),
    .VSS(VGND),
    .A1(_1865_),
    .A2(_1888_));
 sg13g2_o21ai_1 _5106_ (.B1(_1861_),
    .VDD(VPWR),
    .Y(_1902_),
    .VSS(VGND),
    .A1(_1819_),
    .A2(_1859_));
 sg13g2_o21ai_1 _5107_ (.B1(_1870_),
    .VDD(VPWR),
    .Y(_1903_),
    .VSS(VGND),
    .A1(_1867_),
    .A2(_1871_));
 sg13g2_nand2_1 _5108_ (.Y(_1904_),
    .A(net852),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5109_ (.Y(_1905_),
    .A(net848),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5110_ (.Y(_1906_),
    .A(net848),
    .B(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5111_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1907_),
    .B(_1905_),
    .A(_1859_));
 sg13g2_xnor2_1 _5112_ (.Y(_1908_),
    .A(_1858_),
    .B(_1906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5113_ (.B(_1908_),
    .A(_1904_),
    .X(_1909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5114_ (.Y(_1910_),
    .A(_1903_),
    .B(_1909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5115_ (.A(_1910_),
    .B_N(_1902_),
    .Y(_1911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5116_ (.B(_1910_),
    .A(_1902_),
    .X(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5117_ (.B1(_1882_),
    .VDD(VPWR),
    .Y(_1913_),
    .VSS(VGND),
    .A1(_1873_),
    .A2(_1883_));
 sg13g2_nand2_1 _5118_ (.Y(_1914_),
    .A(net846),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5119_ (.Y(_1915_),
    .A(net787),
    .B(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5120_ (.Y(_1916_),
    .A(net789),
    .B(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5121_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1917_),
    .B(_1915_),
    .A(_1869_));
 sg13g2_and2_1 _5122_ (.A(_1868_),
    .B(_1916_),
    .X(_1918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5123_ (.Y(_1919_),
    .A(_1868_),
    .B(_1916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5124_ (.Y(_1920_),
    .A(_1914_),
    .B(_1919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5125_ (.B1(_1877_),
    .VDD(VPWR),
    .Y(_1921_),
    .VSS(VGND),
    .A1(_1875_),
    .A2(_1878_));
 sg13g2_nand2_1 _5126_ (.Y(_1922_),
    .A(net791),
    .B(net998),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5127_ (.A(net794),
    .B(net791),
    .C(net839),
    .D(net997),
    .X(_1923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5128_ (.Y(_1924_),
    .B1(net998),
    .B2(net793),
    .A2(net838),
    .A1(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5129_ (.A(_1923_),
    .B(_1924_),
    .Y(_1925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5130_ (.Y(_1926_),
    .A(_1921_),
    .B(_1925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5131_ (.Y(_1927_),
    .A(_1921_),
    .B(_1925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5132_ (.B(_1927_),
    .A(_1920_),
    .X(_1928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5133_ (.Y(_1929_),
    .A(_1913_),
    .B(_1928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5134_ (.Y(_1930_),
    .A(_1913_),
    .B(_1928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5135_ (.B(_1930_),
    .A(_1912_),
    .X(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5136_ (.Y(_1932_),
    .A(_1901_),
    .B(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5137_ (.Y(_1933_),
    .A(_1901_),
    .B(_1931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5138_ (.Y(_1934_),
    .B(_1900_),
    .A_N(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5139_ (.B(_1933_),
    .A(_1900_),
    .X(_1935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1891_),
    .A2(_1894_),
    .Y(_1936_),
    .B1(_1935_));
 sg13g2_a21o_1 _5141_ (.A2(_1894_),
    .A1(_1891_),
    .B1(_1935_),
    .X(_1937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _5142_ (.X(_1938_),
    .A(_1891_),
    .B(_1894_),
    .C(_1935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5143_ (.A(_1936_),
    .B(_1938_),
    .Y(_1939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5144_ (.Y(_1940_),
    .A(_1896_),
    .B(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5145_ (.B(_1940_),
    .A(_1939_),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5146_ (.A2(_1909_),
    .A1(_1903_),
    .B1(_1911_),
    .X(_1941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5147_ (.B1(_1929_),
    .VDD(VPWR),
    .Y(_1942_),
    .VSS(VGND),
    .A1(_1912_),
    .A2(_1930_));
 sg13g2_o21ai_1 _5148_ (.B1(_1907_),
    .VDD(VPWR),
    .Y(_1943_),
    .VSS(VGND),
    .A1(_1904_),
    .A2(_1908_));
 sg13g2_o21ai_1 _5149_ (.B1(_1917_),
    .VDD(VPWR),
    .Y(_1944_),
    .VSS(VGND),
    .A1(_1914_),
    .A2(_1918_));
 sg13g2_nand2_1 _5150_ (.Y(_1945_),
    .A(net850),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5151_ (.Y(_1946_),
    .A(net846),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5152_ (.Y(_1947_),
    .A(net846),
    .B(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5153_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1948_),
    .B(_1946_),
    .A(_1906_));
 sg13g2_xnor2_1 _5154_ (.Y(_1949_),
    .A(_1905_),
    .B(_1947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5155_ (.B(_1949_),
    .A(_1945_),
    .X(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5156_ (.Y(_1951_),
    .A(_1944_),
    .B(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5157_ (.A(_1951_),
    .B_N(_1943_),
    .Y(_1952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5158_ (.B(_1951_),
    .A(_1943_),
    .X(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5159_ (.B1(_1926_),
    .VDD(VPWR),
    .Y(_1954_),
    .VSS(VGND),
    .A1(_1920_),
    .A2(_1927_));
 sg13g2_a21oi_1 _5160_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net794),
    .A2(net838),
    .Y(_1955_),
    .B1(_1922_));
 sg13g2_nand2_1 _5161_ (.Y(_1956_),
    .A(net844),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5162_ (.Y(_1957_),
    .A(net787),
    .B(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5163_ (.Y(_1958_),
    .A(net789),
    .B(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5164_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1959_),
    .B(_1957_),
    .A(_1916_));
 sg13g2_xnor2_1 _5165_ (.Y(_1960_),
    .A(_1915_),
    .B(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5166_ (.B(_1960_),
    .A(_1956_),
    .X(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5167_ (.Y(_1962_),
    .A(_1955_),
    .B(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5168_ (.Y(_1963_),
    .B(_1954_),
    .A_N(_1962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5169_ (.B(_1962_),
    .A(_1954_),
    .X(_1964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5170_ (.B(_1964_),
    .A(_1953_),
    .X(_1965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5171_ (.Y(_1966_),
    .A(_1942_),
    .B(_1965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5172_ (.B(_1965_),
    .A(_1942_),
    .X(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5173_ (.Y(_1968_),
    .A(_1941_),
    .B(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5174_ (.Y(_1969_),
    .A(_1941_),
    .B(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5175_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1932_),
    .A2(_1934_),
    .Y(_1970_),
    .B1(_1969_));
 sg13g2_nand3_1 _5176_ (.B(_1934_),
    .C(_1969_),
    .A(_1932_),
    .Y(_1971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5177_ (.A(_1970_),
    .B_N(_1971_),
    .Y(_1972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5178_ (.B(_1853_),
    .C(_1898_),
    .A(_1852_),
    .Y(_1973_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1939_));
 sg13g2_a21oi_1 _5179_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1896_),
    .A2(_1937_),
    .Y(_1974_),
    .B1(_1938_));
 sg13g2_nand2b_1 _5180_ (.Y(_1975_),
    .B(_1973_),
    .A_N(_1974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5181_ (.B(_1975_),
    .A(_1972_),
    .X(_0150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5182_ (.A2(_1950_),
    .A1(_1944_),
    .B1(_1952_),
    .X(_1976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5183_ (.B1(_1963_),
    .VDD(VPWR),
    .Y(_1977_),
    .VSS(VGND),
    .A1(_1953_),
    .A2(_1964_));
 sg13g2_a21o_1 _5184_ (.A2(_1961_),
    .A1(_1955_),
    .B1(_1923_),
    .X(_1978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5185_ (.Y(_1979_),
    .A(net785),
    .B(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5186_ (.Y(_1980_),
    .A(net789),
    .B(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5187_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1981_),
    .B(_1980_),
    .A(_1957_));
 sg13g2_xnor2_1 _5188_ (.Y(_1982_),
    .A(_1957_),
    .B(_1980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5189_ (.B(_1982_),
    .A(_1979_),
    .X(_1983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5190_ (.Y(_1984_),
    .A(_1978_),
    .B(_1983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5191_ (.B1(_1948_),
    .VDD(VPWR),
    .Y(_1985_),
    .VSS(VGND),
    .A1(_1945_),
    .A2(_1949_));
 sg13g2_inv_1 _5192_ (.VDD(VPWR),
    .Y(_1986_),
    .A(_1985_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5193_ (.B1(_1959_),
    .VDD(VPWR),
    .Y(_1987_),
    .VSS(VGND),
    .A1(_1956_),
    .A2(_1960_));
 sg13g2_nand2_1 _5194_ (.Y(_1988_),
    .A(net848),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5195_ (.Y(_1989_),
    .A(net844),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5196_ (.Y(_1990_),
    .A(net844),
    .B(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5197_ (.B(_1990_),
    .A(_1946_),
    .X(_1991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5198_ (.Y(_1992_),
    .B(_1991_),
    .A_N(_1988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5199_ (.Y(_1993_),
    .A(_1988_),
    .B(_1991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5200_ (.Y(_1994_),
    .A(_1987_),
    .B(_1993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5201_ (.Y(_1995_),
    .A(_1987_),
    .B(_1993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5202_ (.Y(_1996_),
    .A(_1986_),
    .B(_1995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5203_ (.A(_1984_),
    .B(_1996_),
    .Y(_1997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5204_ (.B(_1996_),
    .A(_1984_),
    .X(_1998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5205_ (.Y(_1999_),
    .A(_1977_),
    .B(_1998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5206_ (.A(_1999_),
    .B_N(_1976_),
    .Y(_2000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5207_ (.B(_1999_),
    .A(_1976_),
    .X(_2001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5208_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1966_),
    .A2(_1968_),
    .Y(_2002_),
    .B1(_2001_));
 sg13g2_nand3_1 _5209_ (.B(_1968_),
    .C(_2001_),
    .A(_1966_),
    .Y(_2003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5210_ (.A(_2002_),
    .B_N(_2003_),
    .Y(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5211_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1972_),
    .A2(_1975_),
    .Y(_2005_),
    .B1(_1970_));
 sg13g2_xnor2_1 _5212_ (.Y(_0151_),
    .A(_2004_),
    .B(_2005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5213_ (.B1(_1994_),
    .VDD(VPWR),
    .Y(_2006_),
    .VSS(VGND),
    .A1(_1986_),
    .A2(_1995_));
 sg13g2_a22oi_1 _5214_ (.Y(_2007_),
    .B1(net997),
    .B2(net787),
    .A2(net838),
    .A1(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5215_ (.Y(_2008_),
    .A(net785),
    .B(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5216_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2009_),
    .B(_2008_),
    .A(_1957_));
 sg13g2_nand2b_1 _5217_ (.Y(_2010_),
    .B(_2009_),
    .A_N(_2007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5218_ (.B1(_1992_),
    .VDD(VPWR),
    .Y(_2011_),
    .VSS(VGND),
    .A1(_1946_),
    .A2(_1990_));
 sg13g2_o21ai_1 _5219_ (.B1(_1981_),
    .VDD(VPWR),
    .Y(_2012_),
    .VSS(VGND),
    .A1(_1979_),
    .A2(_1982_));
 sg13g2_nand2_1 _5220_ (.Y(_2013_),
    .A(net846),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5221_ (.Y(_2014_),
    .A(net841),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5222_ (.Y(_2015_),
    .A(net841),
    .B(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5223_ (.B(_2015_),
    .A(_1989_),
    .X(_2016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5224_ (.Y(_2017_),
    .B(_2016_),
    .A_N(_2013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5225_ (.Y(_2018_),
    .A(_2013_),
    .B(_2016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5226_ (.Y(_2019_),
    .A(_2012_),
    .B(_2018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5227_ (.A(_2019_),
    .B_N(_2011_),
    .Y(_2020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5228_ (.B(_2019_),
    .A(_2011_),
    .X(_2021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5229_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2022_),
    .B(_2021_),
    .A(_2010_));
 sg13g2_xor2_1 _5230_ (.B(_2021_),
    .A(_2010_),
    .X(_2023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5231_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1978_),
    .A2(_1983_),
    .Y(_2024_),
    .B1(_1997_));
 sg13g2_nor2b_1 _5232_ (.A(_2024_),
    .B_N(_2023_),
    .Y(_2025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5233_ (.Y(_2026_),
    .A(_2023_),
    .B(_2024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5234_ (.Y(_2027_),
    .A(_2006_),
    .B(_2026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5235_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1977_),
    .A2(_1998_),
    .Y(_2028_),
    .B1(_2000_));
 sg13g2_nor2_1 _5236_ (.A(_2027_),
    .B(_2028_),
    .Y(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5237_ (.B(_2028_),
    .A(_2027_),
    .X(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5238_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1970_),
    .A2(_2003_),
    .Y(_2031_),
    .B1(_2002_));
 sg13g2_nor2b_1 _5239_ (.A(_1974_),
    .B_N(_2031_),
    .Y(_2032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5240_ (.B1(_2003_),
    .VDD(VPWR),
    .Y(_2033_),
    .VSS(VGND),
    .A1(_1971_),
    .A2(_2002_));
 sg13g2_a21oi_2 _5241_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2033_),
    .Y(_2034_),
    .A2(_2032_),
    .A1(_1973_));
 sg13g2_xor2_1 _5242_ (.B(_2034_),
    .A(_2030_),
    .X(_0152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5243_ (.A2(_2026_),
    .A1(_2006_),
    .B1(_2025_),
    .X(_2035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5244_ (.A2(_2018_),
    .A1(_2012_),
    .B1(_2020_),
    .X(_2036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5245_ (.B1(_2017_),
    .VDD(VPWR),
    .Y(_2037_),
    .VSS(VGND),
    .A1(_1989_),
    .A2(_2015_));
 sg13g2_nand2_1 _5246_ (.Y(_2038_),
    .A(net844),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5247_ (.Y(_2039_),
    .A(net838),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5248_ (.Y(_2040_),
    .A(net783),
    .B(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5249_ (.B(_2040_),
    .A(_2014_),
    .X(_2041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5250_ (.Y(_2042_),
    .B(_2041_),
    .A_N(_2038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5251_ (.Y(_2043_),
    .A(_2038_),
    .B(_2041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5252_ (.A(_2009_),
    .B_N(_2043_),
    .Y(_2044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5253_ (.Y(_2045_),
    .A(_2009_),
    .B(_2043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5254_ (.Y(_2046_),
    .A(_2037_),
    .B(_2045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5255_ (.A(_2008_),
    .B(_2046_),
    .Y(_2047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5256_ (.B(_2046_),
    .A(_2008_),
    .X(_2048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5257_ (.Y(_2049_),
    .B(_2048_),
    .A_N(_2022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5258_ (.Y(_2050_),
    .A(_2022_),
    .B(_2048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5259_ (.Y(_2051_),
    .A(_2036_),
    .B(_2050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5260_ (.Y(_2052_),
    .A(_2036_),
    .B(_2050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5261_ (.A(_2052_),
    .B_N(_2035_),
    .Y(_2053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5262_ (.Y(_2054_),
    .B(_2052_),
    .A_N(_2035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5263_ (.A(_2053_),
    .B_N(_2054_),
    .Y(_2055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5264_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2030_),
    .A2(_2034_),
    .Y(_2056_),
    .B1(_2029_));
 sg13g2_xnor2_1 _5265_ (.Y(_0153_),
    .A(_2055_),
    .B(_2056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5266_ (.A(_2030_),
    .B(_2055_),
    .X(_2057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5267_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2034_),
    .C1(_2053_),
    .B1(_2057_),
    .A1(_2029_),
    .Y(_2058_),
    .A2(_2054_));
 sg13g2_and2_1 _5268_ (.A(_2049_),
    .B(_2051_),
    .X(_2059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5269_ (.A2(_2045_),
    .A1(_2037_),
    .B1(_2044_),
    .X(_2060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5270_ (.Y(_2061_),
    .A(net841),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5271_ (.Y(_2062_),
    .A(net782),
    .B(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5272_ (.Y(_2063_),
    .A(net783),
    .B(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5273_ (.B(_2063_),
    .A(_2039_),
    .X(_2064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5274_ (.Y(_2065_),
    .B(_2064_),
    .A_N(_2061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5275_ (.Y(_2066_),
    .A(_2061_),
    .B(_2064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5276_ (.B1(_2042_),
    .VDD(VPWR),
    .Y(_2067_),
    .VSS(VGND),
    .A1(_2014_),
    .A2(_2040_));
 sg13g2_nand2_1 _5277_ (.Y(_2068_),
    .A(_2066_),
    .B(_2067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5278_ (.B(_2067_),
    .A(_2066_),
    .X(_2069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5279_ (.Y(_2070_),
    .A(_2047_),
    .B(_2069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5280_ (.A(_2070_),
    .B_N(_2060_),
    .Y(_2071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5281_ (.B(_2070_),
    .A(_2060_),
    .X(_2072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5282_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2073_),
    .B(_2072_),
    .A(_2059_));
 sg13g2_xor2_1 _5283_ (.B(_2072_),
    .A(_2059_),
    .X(_2074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5284_ (.VDD(VPWR),
    .Y(_2075_),
    .A(_2074_),
    .VSS(VGND));
 sg13g2_xnor2_1 _5285_ (.Y(_0154_),
    .A(_2058_),
    .B(_2074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5286_ (.B1(_2073_),
    .VDD(VPWR),
    .Y(_2076_),
    .VSS(VGND),
    .A1(_2058_),
    .A2(_2075_));
 sg13g2_a21oi_1 _5287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2047_),
    .A2(_2069_),
    .Y(_2077_),
    .B1(_2071_));
 sg13g2_o21ai_1 _5288_ (.B1(_2065_),
    .VDD(VPWR),
    .Y(_2078_),
    .VSS(VGND),
    .A1(_2039_),
    .A2(_2063_));
 sg13g2_nand2_1 _5289_ (.Y(_2079_),
    .A(net838),
    .B(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5290_ (.B(_2079_),
    .A(_2062_),
    .X(_2080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5291_ (.Y(_2081_),
    .A(_2078_),
    .B(_2080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5292_ (.Y(_2082_),
    .A(_2068_),
    .B(_2081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5293_ (.Y(_2083_),
    .A(_2077_),
    .B(_2082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5294_ (.Y(_0155_),
    .A(_2076_),
    .B(_2083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5295_ (.Y(_2084_),
    .A(\mac1.sum_lvl2_ff[19] ),
    .B(net265),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5296_ (.Y(_2085_),
    .A(\mac1.sum_lvl2_ff[20] ),
    .B(net332),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5297_ (.A(\mac1.sum_lvl2_ff[20] ),
    .B(net332),
    .Y(_2086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5298_ (.B(net332),
    .A(\mac1.sum_lvl2_ff[20] ),
    .X(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5299_ (.Y(_0007_),
    .A(_2084_),
    .B(net333),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5300_ (.B1(_2085_),
    .VDD(VPWR),
    .Y(_2088_),
    .VSS(VGND),
    .A1(_2084_),
    .A2(_2086_));
 sg13g2_and2_1 _5301_ (.A(\mac1.sum_lvl2_ff[21] ),
    .B(net415),
    .X(_2089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5302_ (.B(net415),
    .A(\mac1.sum_lvl2_ff[21] ),
    .X(_2090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5303_ (.B(net416),
    .A(_2088_),
    .X(_0008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5304_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2088_),
    .A2(_2090_),
    .Y(_2091_),
    .B1(_2089_));
 sg13g2_nand2_1 _5305_ (.Y(_2092_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(\mac1.sum_lvl2_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5306_ (.Y(_2093_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5307_ (.B(net495),
    .A(_2091_),
    .X(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5308_ (.B1(_2092_),
    .VDD(VPWR),
    .Y(_2094_),
    .VSS(VGND),
    .A1(_2091_),
    .A2(_2093_));
 sg13g2_and2_1 _5309_ (.A(\mac1.sum_lvl2_ff[23] ),
    .B(\mac1.sum_lvl2_ff[4] ),
    .X(_2095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5310_ (.B(net533),
    .A(\mac1.sum_lvl2_ff[23] ),
    .X(_2096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5311_ (.B(net534),
    .A(_2094_),
    .X(_0010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5312_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2094_),
    .A2(_2096_),
    .Y(_2097_),
    .B1(_2095_));
 sg13g2_nor2_1 _5313_ (.A(\mac1.sum_lvl2_ff[24] ),
    .B(\mac1.sum_lvl2_ff[5] ),
    .Y(_2098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5314_ (.B(net529),
    .A(\mac1.sum_lvl2_ff[24] ),
    .X(_2099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5315_ (.Y(_0011_),
    .A(_2097_),
    .B(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5316_ (.A(\mac1.sum_lvl2_ff[25] ),
    .B(\mac1.sum_lvl2_ff[6] ),
    .X(_2100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5317_ (.Y(_2101_),
    .A(\mac1.sum_lvl2_ff[25] ),
    .B(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5318_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2096_),
    .C1(_2095_),
    .B1(_2094_),
    .A1(\mac1.sum_lvl2_ff[24] ),
    .Y(_2102_),
    .A2(\mac1.sum_lvl2_ff[5] ));
 sg13g2_nor3_1 _5319_ (.A(_2098_),
    .B(_2101_),
    .C(_2102_),
    .Y(_2103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5320_ (.B1(net515),
    .VDD(VPWR),
    .Y(_2104_),
    .VSS(VGND),
    .A1(_2098_),
    .A2(_2102_));
 sg13g2_nor2b_2 _5321_ (.A(_2103_),
    .B_N(net516),
    .Y(_0012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5322_ (.Y(_2105_),
    .A(net499),
    .B(\mac1.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5323_ (.B(\mac1.sum_lvl2_ff[7] ),
    .A(\mac1.sum_lvl2_ff[26] ),
    .X(_2106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5324_ (.B1(_2106_),
    .VDD(VPWR),
    .Y(_2107_),
    .VSS(VGND),
    .A1(_2100_),
    .A2(_2103_));
 sg13g2_or3_1 _5325_ (.A(_2100_),
    .B(_2103_),
    .C(_2106_),
    .X(_2108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5326_ (.A(_2107_),
    .B(_2108_),
    .X(_0013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5327_ (.Y(_2109_),
    .A(\mac1.sum_lvl2_ff[27] ),
    .B(\mac1.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5328_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2105_),
    .A2(_2107_),
    .Y(_2110_),
    .B1(_2109_));
 sg13g2_nand3_1 _5329_ (.B(_2107_),
    .C(_2109_),
    .A(net500),
    .Y(_2111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _5330_ (.A(_2110_),
    .B_N(_2111_),
    .Y(_0014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5331_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.sum_lvl2_ff[27] ),
    .A2(\mac1.sum_lvl2_ff[8] ),
    .Y(_2112_),
    .B1(_2110_));
 sg13g2_nor2_1 _5332_ (.A(\mac1.sum_lvl2_ff[28] ),
    .B(\mac1.sum_lvl2_ff[9] ),
    .Y(_2113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5333_ (.B(net546),
    .A(\mac1.sum_lvl2_ff[28] ),
    .X(_2114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5334_ (.Y(_0015_),
    .A(_2112_),
    .B(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5335_ (.A(\mac1.sum_lvl2_ff[29] ),
    .B(net548),
    .X(_2115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5336_ (.B(net537),
    .A(\mac1.sum_lvl2_ff[29] ),
    .X(_2116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5337_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mac1.sum_lvl2_ff[9] ),
    .C1(_2110_),
    .B1(\mac1.sum_lvl2_ff[28] ),
    .A1(\mac1.sum_lvl2_ff[27] ),
    .Y(_2117_),
    .A2(\mac1.sum_lvl2_ff[8] ));
 sg13g2_nor2_1 _5338_ (.A(_2113_),
    .B(_2117_),
    .Y(_2118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5339_ (.B(_2118_),
    .A(net538),
    .X(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5340_ (.A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ),
    .X(_2119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5341_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2120_),
    .B(\mac1.sum_lvl2_ff[11] ),
    .A(\mac1.sum_lvl2_ff[30] ));
 sg13g2_nor2b_1 _5342_ (.A(_2119_),
    .B_N(_2120_),
    .Y(_2121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5343_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2116_),
    .A2(_2118_),
    .Y(_2122_),
    .B1(_2115_));
 sg13g2_xnor2_1 _5344_ (.Y(_0002_),
    .A(_2121_),
    .B(_2122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5345_ (.Y(_2123_),
    .A(_2116_),
    .B(_2121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5346_ (.A(_2113_),
    .B(_2117_),
    .C(_2123_),
    .Y(_2124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5347_ (.A2(_2120_),
    .A1(_2115_),
    .B1(_2119_),
    .X(_2125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5348_ (.A(_2124_),
    .B(_2125_),
    .Y(_2126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5349_ (.Y(_2127_),
    .A(\mac1.sum_lvl2_ff[31] ),
    .B(\mac1.sum_lvl2_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5350_ (.B(net535),
    .A(\mac1.sum_lvl2_ff[31] ),
    .X(_2128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5351_ (.B1(_2128_),
    .VDD(VPWR),
    .Y(_2129_),
    .VSS(VGND),
    .A1(_2124_),
    .A2(_2125_));
 sg13g2_xnor2_1 _5352_ (.Y(_0003_),
    .A(_2126_),
    .B(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5353_ (.Y(_2130_),
    .A(\mac1.sum_lvl2_ff[32] ),
    .B(net478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5354_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2127_),
    .A2(_2129_),
    .Y(_2131_),
    .B1(net479));
 sg13g2_nand3_1 _5355_ (.B(_2129_),
    .C(net479),
    .A(_2127_),
    .Y(_2132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _5356_ (.A(net480),
    .B_N(_2132_),
    .Y(_0004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5357_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.sum_lvl2_ff[32] ),
    .A2(\mac1.sum_lvl2_ff[13] ),
    .Y(_2133_),
    .B1(_2131_));
 sg13g2_nand2_1 _5358_ (.Y(_2134_),
    .A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5359_ (.A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .Y(_2135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5360_ (.B(net468),
    .A(\mac1.sum_lvl2_ff[33] ),
    .X(_2136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5361_ (.Y(_0005_),
    .A(_2133_),
    .B(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5362_ (.B1(_2134_),
    .VDD(VPWR),
    .Y(_2137_),
    .VSS(VGND),
    .A1(_2133_),
    .A2(_2135_));
 sg13g2_xnor2_1 _5363_ (.Y(_2138_),
    .A(\mac1.sum_lvl2_ff[34] ),
    .B(net285),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5364_ (.Y(_0006_),
    .A(_2137_),
    .B(net286),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5365_ (.B(net265),
    .A(\mac1.sum_lvl2_ff[19] ),
    .X(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5366_ (.Y(_2139_),
    .A(net429),
    .B(net283),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5367_ (.Y(_2140_),
    .A(\mac1.sum_lvl3_ff[21] ),
    .B(\mac1.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5368_ (.A(\mac1.sum_lvl3_ff[21] ),
    .B(\mac1.sum_lvl3_ff[1] ),
    .Y(_2141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5369_ (.B(\mac1.sum_lvl3_ff[1] ),
    .A(\mac1.sum_lvl3_ff[21] ),
    .X(_2142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5370_ (.Y(_0023_),
    .A(_2139_),
    .B(_2142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5371_ (.B1(_2140_),
    .VDD(VPWR),
    .Y(_2143_),
    .VSS(VGND),
    .A1(_2139_),
    .A2(_2141_));
 sg13g2_and2_1 _5372_ (.A(\mac1.sum_lvl3_ff[22] ),
    .B(\mac1.sum_lvl3_ff[2] ),
    .X(_2144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5373_ (.B(net433),
    .A(\mac1.sum_lvl3_ff[22] ),
    .X(_2145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5374_ (.B(net434),
    .A(_2143_),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _5375_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2144_),
    .Y(_2146_),
    .A2(_2145_),
    .A1(_2143_));
 sg13g2_nand2_1 _5376_ (.Y(_2147_),
    .A(\mac1.sum_lvl3_ff[23] ),
    .B(\mac1.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5377_ (.Y(_2148_),
    .A(\mac1.sum_lvl3_ff[23] ),
    .B(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5378_ (.B(net384),
    .A(_2146_),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5379_ (.B1(_2147_),
    .VDD(VPWR),
    .Y(_2149_),
    .VSS(VGND),
    .A1(_2146_),
    .A2(_2148_));
 sg13g2_and2_1 _5380_ (.A(\mac1.sum_lvl3_ff[24] ),
    .B(\mac1.sum_lvl3_ff[4] ),
    .X(_2150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5381_ (.B(net353),
    .A(\mac1.sum_lvl3_ff[24] ),
    .X(_2151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5382_ (.B(net354),
    .A(_2149_),
    .X(_0026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5383_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2149_),
    .A2(_2151_),
    .Y(_2152_),
    .B1(_2150_));
 sg13g2_nor2_1 _5384_ (.A(\mac1.sum_lvl3_ff[25] ),
    .B(net317),
    .Y(_2153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5385_ (.B(net317),
    .A(\mac1.sum_lvl3_ff[25] ),
    .X(_2154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5386_ (.Y(_0027_),
    .A(_2152_),
    .B(net318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5387_ (.A(\mac1.sum_lvl3_ff[26] ),
    .B(net483),
    .X(_2155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5388_ (.Y(_2156_),
    .A(\mac1.sum_lvl3_ff[26] ),
    .B(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5389_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2151_),
    .C1(_2150_),
    .B1(_2149_),
    .A1(\mac1.sum_lvl3_ff[25] ),
    .Y(_2157_),
    .A2(\mac1.sum_lvl3_ff[5] ));
 sg13g2_nor3_1 _5390_ (.A(_2153_),
    .B(net484),
    .C(_2157_),
    .Y(_2158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5391_ (.B1(net484),
    .VDD(VPWR),
    .Y(_2159_),
    .VSS(VGND),
    .A1(_2153_),
    .A2(_2157_));
 sg13g2_nor2b_1 _5392_ (.A(_2158_),
    .B_N(net485),
    .Y(_0028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5393_ (.Y(_2160_),
    .A(\mac1.sum_lvl3_ff[27] ),
    .B(\mac1.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5394_ (.B(net518),
    .A(\mac1.sum_lvl3_ff[27] ),
    .X(_2161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5395_ (.B1(net519),
    .VDD(VPWR),
    .Y(_2162_),
    .VSS(VGND),
    .A1(_2155_),
    .A2(_2158_));
 sg13g2_or3_1 _5396_ (.A(_2155_),
    .B(_2158_),
    .C(net519),
    .X(_2163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5397_ (.A(net520),
    .B(_2163_),
    .X(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5398_ (.Y(_2164_),
    .A(\mac1.sum_lvl3_ff[28] ),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5399_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2160_),
    .A2(_2162_),
    .Y(_2165_),
    .B1(net406));
 sg13g2_nand3_1 _5400_ (.B(_2162_),
    .C(net406),
    .A(_2160_),
    .Y(_2166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5401_ (.A(net407),
    .B_N(_2166_),
    .Y(_0030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5402_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.sum_lvl3_ff[28] ),
    .A2(\mac1.sum_lvl3_ff[8] ),
    .Y(_2167_),
    .B1(_2165_));
 sg13g2_nand2_1 _5403_ (.Y(_2168_),
    .A(\mac1.sum_lvl3_ff[29] ),
    .B(net293),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5404_ (.A(\mac1.sum_lvl3_ff[29] ),
    .B(net293),
    .Y(_2169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5405_ (.B(net293),
    .A(\mac1.sum_lvl3_ff[29] ),
    .X(_2170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5406_ (.Y(_0031_),
    .A(_2167_),
    .B(net294),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5407_ (.B1(_2168_),
    .VDD(VPWR),
    .Y(_2171_),
    .VSS(VGND),
    .A1(_2167_),
    .A2(_2169_));
 sg13g2_nand2_1 _5408_ (.Y(_2172_),
    .A(\mac1.sum_lvl3_ff[30] ),
    .B(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5409_ (.Y(_2173_),
    .A(\mac1.sum_lvl3_ff[30] ),
    .B(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5410_ (.Y(_2174_),
    .B(_2171_),
    .A_N(_2173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5411_ (.Y(_0017_),
    .A(_2171_),
    .B(net378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5412_ (.A(\mac1.sum_lvl3_ff[31] ),
    .B(\mac1.sum_lvl3_ff[11] ),
    .Y(_2175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5413_ (.Y(_2176_),
    .A(\mac1.sum_lvl3_ff[31] ),
    .B(net393),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5414_ (.Y(_2177_),
    .A(_2172_),
    .B(_2174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5415_ (.Y(_0018_),
    .A(net394),
    .B(_2177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5416_ (.A(_2173_),
    .B(_2176_),
    .Y(_2178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5417_ (.A(_2172_),
    .B(_2175_),
    .Y(_2179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5418_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2178_),
    .C1(_2179_),
    .B1(_2171_),
    .A1(\mac1.sum_lvl3_ff[31] ),
    .Y(_2180_),
    .A2(\mac1.sum_lvl3_ff[11] ));
 sg13g2_nand2_1 _5419_ (.Y(_2181_),
    .A(\mac1.sum_lvl3_ff[32] ),
    .B(net323),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5420_ (.A(\mac1.sum_lvl3_ff[32] ),
    .B(net323),
    .Y(_2182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5421_ (.B(net323),
    .A(\mac1.sum_lvl3_ff[32] ),
    .X(_2183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5422_ (.Y(_0019_),
    .A(_2180_),
    .B(net324),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5423_ (.B1(_2181_),
    .VDD(VPWR),
    .Y(_2184_),
    .VSS(VGND),
    .A1(_2180_),
    .A2(_2182_));
 sg13g2_or2_1 _5424_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2185_),
    .B(net341),
    .A(\mac1.sum_lvl3_ff[33] ));
 sg13g2_and2_1 _5425_ (.A(\mac1.sum_lvl3_ff[33] ),
    .B(net341),
    .X(_2186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5426_ (.Y(_2187_),
    .A(\mac1.sum_lvl3_ff[33] ),
    .B(net341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5427_ (.Y(_0020_),
    .A(_2184_),
    .B(net342),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5428_ (.Y(_2188_),
    .A(\mac1.sum_lvl3_ff[34] ),
    .B(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5429_ (.A(\mac1.sum_lvl3_ff[34] ),
    .B(net373),
    .Y(_2189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5430_ (.B(net373),
    .A(\mac1.sum_lvl3_ff[34] ),
    .X(_2190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5431_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2184_),
    .A2(_2185_),
    .Y(_2191_),
    .B1(_2186_));
 sg13g2_xnor2_1 _5432_ (.Y(_0021_),
    .A(net374),
    .B(_2191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5433_ (.B1(_2188_),
    .VDD(VPWR),
    .Y(_2192_),
    .VSS(VGND),
    .A1(_2189_),
    .A2(_2191_));
 sg13g2_xnor2_1 _5434_ (.Y(_2193_),
    .A(net409),
    .B(\mac1.sum_lvl3_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5435_ (.Y(_0022_),
    .A(_2192_),
    .B(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5436_ (.B(net283),
    .A(\mac1.sum_lvl3_ff[20] ),
    .X(_0016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5437_ (.Y(_2194_),
    .A(net291),
    .B(net267),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5438_ (.Y(_2195_),
    .A(\mac2.sum_lvl2_ff[20] ),
    .B(\mac2.sum_lvl2_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5439_ (.A(\mac2.sum_lvl2_ff[20] ),
    .B(\mac2.sum_lvl2_ff[1] ),
    .Y(_2196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5440_ (.B(\mac2.sum_lvl2_ff[1] ),
    .A(\mac2.sum_lvl2_ff[20] ),
    .X(_2197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5441_ (.Y(_0039_),
    .A(_2194_),
    .B(_2197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5442_ (.B1(_2195_),
    .VDD(VPWR),
    .Y(_2198_),
    .VSS(VGND),
    .A1(_2194_),
    .A2(_2196_));
 sg13g2_and2_1 _5443_ (.A(\mac2.sum_lvl2_ff[21] ),
    .B(net320),
    .X(_2199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5444_ (.B(net320),
    .A(\mac2.sum_lvl2_ff[21] ),
    .X(_2200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5445_ (.B(net321),
    .A(_2198_),
    .X(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5446_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2198_),
    .A2(net321),
    .Y(_2201_),
    .B1(_2199_));
 sg13g2_nand2_1 _5447_ (.Y(_2202_),
    .A(\mac2.sum_lvl2_ff[22] ),
    .B(net360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5448_ (.Y(_2203_),
    .A(\mac2.sum_lvl2_ff[22] ),
    .B(net360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5449_ (.B(net361),
    .A(_2201_),
    .X(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5450_ (.B1(_2202_),
    .VDD(VPWR),
    .Y(_2204_),
    .VSS(VGND),
    .A1(_2201_),
    .A2(_2203_));
 sg13g2_and2_1 _5451_ (.A(\mac2.sum_lvl2_ff[23] ),
    .B(\mac2.sum_lvl2_ff[4] ),
    .X(_2205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5452_ (.B(net461),
    .A(\mac2.sum_lvl2_ff[23] ),
    .X(_2206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5453_ (.B(net462),
    .A(_2204_),
    .X(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5454_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2204_),
    .A2(_2206_),
    .Y(_2207_),
    .B1(_2205_));
 sg13g2_nor2_1 _5455_ (.A(\mac2.sum_lvl2_ff[24] ),
    .B(net448),
    .Y(_2208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5456_ (.B(net448),
    .A(\mac2.sum_lvl2_ff[24] ),
    .X(_2209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5457_ (.Y(_0043_),
    .A(_2207_),
    .B(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5458_ (.A(\mac2.sum_lvl2_ff[25] ),
    .B(\mac2.sum_lvl2_ff[6] ),
    .X(_2210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5459_ (.Y(_2211_),
    .A(\mac2.sum_lvl2_ff[25] ),
    .B(net524),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5460_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2206_),
    .C1(_2205_),
    .B1(_2204_),
    .A1(\mac2.sum_lvl2_ff[24] ),
    .Y(_2212_),
    .A2(\mac2.sum_lvl2_ff[5] ));
 sg13g2_nor3_2 _5461_ (.A(_2208_),
    .B(net525),
    .C(_2212_),
    .Y(_2213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5462_ (.B1(net525),
    .VDD(VPWR),
    .Y(_2214_),
    .VSS(VGND),
    .A1(_2208_),
    .A2(_2212_));
 sg13g2_nor2b_2 _5463_ (.A(_2213_),
    .B_N(net526),
    .Y(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5464_ (.Y(_2215_),
    .A(\mac2.sum_lvl2_ff[26] ),
    .B(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5465_ (.B(\mac2.sum_lvl2_ff[7] ),
    .A(\mac2.sum_lvl2_ff[26] ),
    .X(_2216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5466_ (.B1(_2216_),
    .VDD(VPWR),
    .Y(_2217_),
    .VSS(VGND),
    .A1(_2210_),
    .A2(_2213_));
 sg13g2_or3_1 _5467_ (.A(_2210_),
    .B(_2213_),
    .C(_2216_),
    .X(_2218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5468_ (.A(_2217_),
    .B(_2218_),
    .X(_0045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5469_ (.Y(_2219_),
    .A(\mac2.sum_lvl2_ff[27] ),
    .B(\mac2.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _5470_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2219_),
    .Y(_2220_),
    .A2(_2217_),
    .A1(net507));
 sg13g2_nand3_1 _5471_ (.B(_2217_),
    .C(_2219_),
    .A(net507),
    .Y(_2221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _5472_ (.A(_2220_),
    .B_N(_2221_),
    .Y(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5473_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac2.sum_lvl2_ff[27] ),
    .A2(\mac2.sum_lvl2_ff[8] ),
    .Y(_2222_),
    .B1(_2220_));
 sg13g2_nor2_1 _5474_ (.A(\mac2.sum_lvl2_ff[28] ),
    .B(\mac2.sum_lvl2_ff[9] ),
    .Y(_2223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5475_ (.B(net542),
    .A(\mac2.sum_lvl2_ff[28] ),
    .X(_2224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5476_ (.Y(_0047_),
    .A(_2222_),
    .B(net543),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5477_ (.A(\mac2.sum_lvl2_ff[29] ),
    .B(\mac2.sum_lvl2_ff[10] ),
    .X(_2225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5478_ (.B(net544),
    .A(\mac2.sum_lvl2_ff[29] ),
    .X(_2226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5479_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mac2.sum_lvl2_ff[9] ),
    .C1(_2220_),
    .B1(\mac2.sum_lvl2_ff[28] ),
    .A1(\mac2.sum_lvl2_ff[27] ),
    .Y(_2227_),
    .A2(\mac2.sum_lvl2_ff[8] ));
 sg13g2_nor2_1 _5480_ (.A(_2223_),
    .B(_2227_),
    .Y(_2228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5481_ (.B(_2228_),
    .A(net545),
    .X(_0033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5482_ (.A(\mac2.sum_lvl2_ff[30] ),
    .B(\mac2.sum_lvl2_ff[11] ),
    .X(_2229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5483_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2230_),
    .B(\mac2.sum_lvl2_ff[11] ),
    .A(\mac2.sum_lvl2_ff[30] ));
 sg13g2_nor2b_1 _5484_ (.A(_2229_),
    .B_N(_2230_),
    .Y(_2231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5485_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2226_),
    .A2(_2228_),
    .Y(_2232_),
    .B1(_2225_));
 sg13g2_xnor2_1 _5486_ (.Y(_0034_),
    .A(_2231_),
    .B(_2232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5487_ (.Y(_2233_),
    .A(_2226_),
    .B(_2231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5488_ (.A(_2223_),
    .B(_2227_),
    .C(_2233_),
    .Y(_2234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5489_ (.A2(_2230_),
    .A1(_2225_),
    .B1(_2229_),
    .X(_2235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5490_ (.A(_2234_),
    .B(_2235_),
    .Y(_2236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5491_ (.Y(_2237_),
    .A(net511),
    .B(\mac2.sum_lvl2_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5492_ (.B(\mac2.sum_lvl2_ff[12] ),
    .A(\mac2.sum_lvl2_ff[31] ),
    .X(_2238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5493_ (.B1(_2238_),
    .VDD(VPWR),
    .Y(_2239_),
    .VSS(VGND),
    .A1(_2234_),
    .A2(_2235_));
 sg13g2_xnor2_1 _5494_ (.Y(_0035_),
    .A(_2236_),
    .B(_2238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5495_ (.Y(_2240_),
    .A(\mac2.sum_lvl2_ff[32] ),
    .B(\mac2.sum_lvl2_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5496_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net512),
    .A2(_2239_),
    .Y(_2241_),
    .B1(_2240_));
 sg13g2_nand3_1 _5497_ (.B(_2239_),
    .C(_2240_),
    .A(net512),
    .Y(_2242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _5498_ (.A(_2241_),
    .B_N(_2242_),
    .Y(_0036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5499_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac2.sum_lvl2_ff[32] ),
    .A2(\mac2.sum_lvl2_ff[13] ),
    .Y(_2243_),
    .B1(_2241_));
 sg13g2_nand2_1 _5500_ (.Y(_2244_),
    .A(\mac2.sum_lvl2_ff[33] ),
    .B(\mac2.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5501_ (.A(\mac2.sum_lvl2_ff[33] ),
    .B(\mac2.sum_lvl2_ff[14] ),
    .Y(_2245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5502_ (.B(\mac2.sum_lvl2_ff[14] ),
    .A(\mac2.sum_lvl2_ff[33] ),
    .X(_2246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5503_ (.Y(_0037_),
    .A(_2243_),
    .B(_2246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5504_ (.B1(_2244_),
    .VDD(VPWR),
    .Y(_2247_),
    .VSS(VGND),
    .A1(_2243_),
    .A2(_2245_));
 sg13g2_xnor2_1 _5505_ (.Y(_2248_),
    .A(\mac2.sum_lvl2_ff[34] ),
    .B(net531),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5506_ (.Y(_0038_),
    .A(_2247_),
    .B(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5507_ (.B(net267),
    .A(\mac2.sum_lvl2_ff[19] ),
    .X(_0032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5508_ (.Y(_2249_),
    .A(net474),
    .B(net305),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5509_ (.Y(_2250_),
    .A(\mac2.sum_lvl3_ff[21] ),
    .B(\mac2.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5510_ (.A(\mac2.sum_lvl3_ff[21] ),
    .B(\mac2.sum_lvl3_ff[1] ),
    .Y(_2251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5511_ (.B(\mac2.sum_lvl3_ff[1] ),
    .A(\mac2.sum_lvl3_ff[21] ),
    .X(_2252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5512_ (.Y(_0055_),
    .A(_2249_),
    .B(_2252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5513_ (.B1(_2250_),
    .VDD(VPWR),
    .Y(_2253_),
    .VSS(VGND),
    .A1(_2249_),
    .A2(_2251_));
 sg13g2_and2_1 _5514_ (.A(\mac2.sum_lvl3_ff[22] ),
    .B(net451),
    .X(_2254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5515_ (.B(net451),
    .A(\mac2.sum_lvl3_ff[22] ),
    .X(_2255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5516_ (.B(net452),
    .A(_2253_),
    .X(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5517_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2253_),
    .A2(_2255_),
    .Y(_2256_),
    .B1(_2254_));
 sg13g2_nand2_1 _5518_ (.Y(_2257_),
    .A(\mac2.sum_lvl3_ff[23] ),
    .B(\mac2.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5519_ (.Y(_2258_),
    .A(\mac2.sum_lvl3_ff[23] ),
    .B(net487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5520_ (.B(net488),
    .A(_2256_),
    .X(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5521_ (.B1(_2257_),
    .VDD(VPWR),
    .Y(_2259_),
    .VSS(VGND),
    .A1(_2256_),
    .A2(_2258_));
 sg13g2_and2_1 _5522_ (.A(\mac2.sum_lvl3_ff[24] ),
    .B(\mac2.sum_lvl3_ff[4] ),
    .X(_2260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5523_ (.B(net454),
    .A(\mac2.sum_lvl3_ff[24] ),
    .X(_2261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5524_ (.B(net455),
    .A(_2259_),
    .X(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5525_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2259_),
    .A2(_2261_),
    .Y(_2262_),
    .B1(_2260_));
 sg13g2_nor2_1 _5526_ (.A(\mac2.sum_lvl3_ff[25] ),
    .B(net418),
    .Y(_2263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5527_ (.B(net418),
    .A(\mac2.sum_lvl3_ff[25] ),
    .X(_2264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5528_ (.Y(_0059_),
    .A(_2262_),
    .B(net419),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5529_ (.A(\mac2.sum_lvl3_ff[26] ),
    .B(\mac2.sum_lvl3_ff[6] ),
    .X(_2265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5530_ (.Y(_2266_),
    .A(\mac2.sum_lvl3_ff[26] ),
    .B(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5531_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2261_),
    .C1(_2260_),
    .B1(_2259_),
    .A1(\mac2.sum_lvl3_ff[25] ),
    .Y(_2267_),
    .A2(net418));
 sg13g2_nor3_1 _5532_ (.A(_2263_),
    .B(net458),
    .C(_2267_),
    .Y(_2268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5533_ (.B1(net458),
    .VDD(VPWR),
    .Y(_2269_),
    .VSS(VGND),
    .A1(_2263_),
    .A2(_2267_));
 sg13g2_nor2b_1 _5534_ (.A(_2268_),
    .B_N(net459),
    .Y(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5535_ (.Y(_2270_),
    .A(net436),
    .B(\mac2.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5536_ (.B(net539),
    .A(net436),
    .X(_2271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5537_ (.B1(_2271_),
    .VDD(VPWR),
    .Y(_2272_),
    .VSS(VGND),
    .A1(_2265_),
    .A2(_2268_));
 sg13g2_or3_1 _5538_ (.A(_2265_),
    .B(_2268_),
    .C(_2271_),
    .X(_2273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5539_ (.A(_2272_),
    .B(net540),
    .X(_0061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5540_ (.Y(_2274_),
    .A(\mac2.sum_lvl3_ff[28] ),
    .B(\mac2.sum_lvl3_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5541_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net437),
    .A2(_2272_),
    .Y(_2275_),
    .B1(_2274_));
 sg13g2_nand3_1 _5542_ (.B(_2272_),
    .C(_2274_),
    .A(net437),
    .Y(_2276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5543_ (.A(_2275_),
    .B_N(net438),
    .Y(_0062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5544_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac2.sum_lvl3_ff[28] ),
    .A2(\mac2.sum_lvl3_ff[8] ),
    .Y(_2277_),
    .B1(_2275_));
 sg13g2_nor2_1 _5545_ (.A(\mac2.sum_lvl3_ff[29] ),
    .B(net338),
    .Y(_2278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5546_ (.B(net338),
    .A(\mac2.sum_lvl3_ff[29] ),
    .X(_2279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5547_ (.Y(_0063_),
    .A(_2277_),
    .B(net339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5548_ (.A(net380),
    .B(\mac2.sum_lvl3_ff[10] ),
    .X(_2280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5549_ (.B(\mac2.sum_lvl3_ff[10] ),
    .A(net380),
    .X(_2281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5550_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net338),
    .C1(_2275_),
    .B1(\mac2.sum_lvl3_ff[29] ),
    .A1(\mac2.sum_lvl3_ff[28] ),
    .Y(_2282_),
    .A2(\mac2.sum_lvl3_ff[8] ));
 sg13g2_nor2_1 _5551_ (.A(_2278_),
    .B(_2282_),
    .Y(_2283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5552_ (.B(_2283_),
    .A(net381),
    .X(_0049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5553_ (.A(net423),
    .B(\mac2.sum_lvl3_ff[11] ),
    .X(_2284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5554_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2285_),
    .B(\mac2.sum_lvl3_ff[11] ),
    .A(net423));
 sg13g2_nor2b_1 _5555_ (.A(net424),
    .B_N(_2285_),
    .Y(_2286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5556_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net381),
    .A2(_2283_),
    .Y(_2287_),
    .B1(_2280_));
 sg13g2_xnor2_1 _5557_ (.Y(_0050_),
    .A(net425),
    .B(_2287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5558_ (.Y(_2288_),
    .A(_2281_),
    .B(_2286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5559_ (.A(_2278_),
    .B(_2282_),
    .C(_2288_),
    .Y(_2289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5560_ (.A2(_2285_),
    .A1(_2280_),
    .B1(_2284_),
    .X(_2290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5561_ (.A(_2289_),
    .B(_2290_),
    .Y(_2291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5562_ (.Y(_2292_),
    .A(\mac2.sum_lvl3_ff[32] ),
    .B(net311),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5563_ (.B(net311),
    .A(\mac2.sum_lvl3_ff[32] ),
    .X(_2293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5564_ (.B1(net312),
    .VDD(VPWR),
    .Y(_2294_),
    .VSS(VGND),
    .A1(_2289_),
    .A2(_2290_));
 sg13g2_xnor2_1 _5565_ (.Y(_0051_),
    .A(_2291_),
    .B(net312),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5566_ (.Y(_2295_),
    .A(\mac2.sum_lvl3_ff[33] ),
    .B(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2292_),
    .A2(_2294_),
    .Y(_2296_),
    .B1(net399));
 sg13g2_nand3_1 _5568_ (.B(_2294_),
    .C(net399),
    .A(_2292_),
    .Y(_2297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5569_ (.A(net400),
    .B_N(_2297_),
    .Y(_0052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5570_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac2.sum_lvl3_ff[33] ),
    .A2(\mac2.sum_lvl3_ff[13] ),
    .Y(_2298_),
    .B1(_2296_));
 sg13g2_nand2_1 _5571_ (.Y(_2299_),
    .A(\mac2.sum_lvl3_ff[34] ),
    .B(net347),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5572_ (.A(\mac2.sum_lvl3_ff[34] ),
    .B(net347),
    .Y(_2300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5573_ (.B(net347),
    .A(\mac2.sum_lvl3_ff[34] ),
    .X(_2301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5574_ (.Y(_0053_),
    .A(_2298_),
    .B(net348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5575_ (.B1(_2299_),
    .VDD(VPWR),
    .Y(_2302_),
    .VSS(VGND),
    .A1(_2298_),
    .A2(_2300_));
 sg13g2_xnor2_1 _5576_ (.Y(_2303_),
    .A(\mac2.sum_lvl3_ff[35] ),
    .B(net367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5577_ (.Y(_0054_),
    .A(_2302_),
    .B(net368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5578_ (.B(net305),
    .A(\mac2.sum_lvl3_ff[20] ),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5579_ (.Y(_2304_),
    .A(\mac1.total_sum[0] ),
    .B(\mac2.total_sum[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5580_ (.Y(_2305_),
    .A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5581_ (.A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .Y(_2306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5582_ (.B(\mac2.total_sum[1] ),
    .A(\mac1.total_sum[1] ),
    .X(_2307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5583_ (.Y(net26),
    .A(_2304_),
    .B(_2307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5584_ (.B1(_2305_),
    .VDD(VPWR),
    .Y(_2308_),
    .VSS(VGND),
    .A1(_2304_),
    .A2(_2306_));
 sg13g2_and2_1 _5585_ (.A(\mac1.total_sum[2] ),
    .B(\mac2.total_sum[2] ),
    .X(_2309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5586_ (.B(\mac2.total_sum[2] ),
    .A(\mac1.total_sum[2] ),
    .X(_2310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5587_ (.B(_2310_),
    .A(_2308_),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5588_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2308_),
    .A2(_2310_),
    .Y(_2311_),
    .B1(_2309_));
 sg13g2_nand2_1 _5589_ (.Y(_2312_),
    .A(\mac1.total_sum[3] ),
    .B(\mac2.total_sum[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5590_ (.Y(_2313_),
    .A(\mac1.total_sum[3] ),
    .B(\mac2.total_sum[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5591_ (.B(_2313_),
    .A(_2311_),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5592_ (.B1(_2312_),
    .VDD(VPWR),
    .Y(_2314_),
    .VSS(VGND),
    .A1(_2311_),
    .A2(_2313_));
 sg13g2_and2_1 _5593_ (.A(\mac1.total_sum[4] ),
    .B(\mac2.total_sum[4] ),
    .X(_2315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5594_ (.B(\mac2.total_sum[4] ),
    .A(\mac1.total_sum[4] ),
    .X(_2316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5595_ (.B(_2316_),
    .A(_2314_),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5596_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2314_),
    .A2(_2316_),
    .Y(_2317_),
    .B1(_2315_));
 sg13g2_nor2_1 _5597_ (.A(\mac1.total_sum[5] ),
    .B(\mac2.total_sum[5] ),
    .Y(_2318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5598_ (.B(\mac2.total_sum[5] ),
    .A(\mac1.total_sum[5] ),
    .X(_2319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5599_ (.Y(net30),
    .A(_2317_),
    .B(_2319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5600_ (.A(\mac1.total_sum[6] ),
    .B(\mac2.total_sum[6] ),
    .X(_2320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5601_ (.Y(_2321_),
    .A(\mac1.total_sum[6] ),
    .B(\mac2.total_sum[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5602_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2316_),
    .C1(_2315_),
    .B1(_2314_),
    .A1(\mac1.total_sum[5] ),
    .Y(_2322_),
    .A2(\mac2.total_sum[5] ));
 sg13g2_nor3_1 _5603_ (.A(_2318_),
    .B(_2321_),
    .C(_2322_),
    .Y(_2323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5604_ (.B1(_2321_),
    .VDD(VPWR),
    .Y(_2324_),
    .VSS(VGND),
    .A1(_2318_),
    .A2(_2322_));
 sg13g2_nor2b_1 _5605_ (.A(_2323_),
    .B_N(_2324_),
    .Y(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5606_ (.Y(_2325_),
    .A(\mac1.total_sum[7] ),
    .B(\mac2.total_sum[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5607_ (.B(\mac2.total_sum[7] ),
    .A(\mac1.total_sum[7] ),
    .X(_2326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5608_ (.B1(_2326_),
    .VDD(VPWR),
    .Y(_2327_),
    .VSS(VGND),
    .A1(_2320_),
    .A2(_2323_));
 sg13g2_or3_1 _5609_ (.A(_2320_),
    .B(_2323_),
    .C(_2326_),
    .X(_2328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5610_ (.A(_2327_),
    .B(_2328_),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5611_ (.Y(_2329_),
    .A(\mac1.total_sum[8] ),
    .B(\mac2.total_sum[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5612_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2325_),
    .A2(_2327_),
    .Y(_2330_),
    .B1(_2329_));
 sg13g2_nand3_1 _5613_ (.B(_2327_),
    .C(_2329_),
    .A(_2325_),
    .Y(_2331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5614_ (.A(_2330_),
    .B_N(_2331_),
    .Y(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5615_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.total_sum[8] ),
    .A2(\mac2.total_sum[8] ),
    .Y(_2332_),
    .B1(_2330_));
 sg13g2_nor2_1 _5616_ (.A(\mac1.total_sum[9] ),
    .B(\mac2.total_sum[9] ),
    .Y(_2333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5617_ (.B(\mac2.total_sum[9] ),
    .A(\mac1.total_sum[9] ),
    .X(_2334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5618_ (.Y(net18),
    .A(_2332_),
    .B(_2334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5619_ (.A(\mac1.total_sum[10] ),
    .B(\mac2.total_sum[10] ),
    .X(_2335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5620_ (.B(\mac2.total_sum[10] ),
    .A(\mac1.total_sum[10] ),
    .X(_2336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5621_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\mac2.total_sum[9] ),
    .C1(_2330_),
    .B1(\mac1.total_sum[9] ),
    .A1(\mac1.total_sum[8] ),
    .Y(_2337_),
    .A2(\mac2.total_sum[8] ));
 sg13g2_nor2_1 _5622_ (.A(_2333_),
    .B(_2337_),
    .Y(_2338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5623_ (.B(_2338_),
    .A(_2336_),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5624_ (.A(\mac1.total_sum[11] ),
    .B(\mac2.total_sum[11] ),
    .X(_2339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5625_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2340_),
    .B(\mac2.total_sum[11] ),
    .A(\mac1.total_sum[11] ));
 sg13g2_nor2b_1 _5626_ (.A(_2339_),
    .B_N(_2340_),
    .Y(_2341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5627_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2336_),
    .A2(_2338_),
    .Y(_2342_),
    .B1(_2335_));
 sg13g2_xnor2_1 _5628_ (.Y(net20),
    .A(_2341_),
    .B(_2342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5629_ (.Y(_2343_),
    .A(_2336_),
    .B(_2341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5630_ (.A(_2333_),
    .B(_2337_),
    .C(_2343_),
    .Y(_2344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5631_ (.A2(_2340_),
    .A1(_2335_),
    .B1(_2339_),
    .X(_2345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5632_ (.A(_2344_),
    .B(_2345_),
    .Y(_2346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5633_ (.Y(_2347_),
    .A(\mac1.total_sum[12] ),
    .B(\mac2.total_sum[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5634_ (.B(\mac2.total_sum[12] ),
    .A(\mac1.total_sum[12] ),
    .X(_2348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5635_ (.B1(_2348_),
    .VDD(VPWR),
    .Y(_2349_),
    .VSS(VGND),
    .A1(_2344_),
    .A2(_2345_));
 sg13g2_xnor2_1 _5636_ (.Y(net21),
    .A(_2346_),
    .B(_2348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5637_ (.Y(_2350_),
    .A(\mac1.total_sum[13] ),
    .B(\mac2.total_sum[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5638_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2347_),
    .A2(_2349_),
    .Y(_2351_),
    .B1(_2350_));
 sg13g2_nand3_1 _5639_ (.B(_2349_),
    .C(_2350_),
    .A(_2347_),
    .Y(_2352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5640_ (.A(_2351_),
    .B_N(_2352_),
    .Y(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.total_sum[13] ),
    .A2(\mac2.total_sum[13] ),
    .Y(_2353_),
    .B1(_2351_));
 sg13g2_nand2_1 _5642_ (.Y(_2354_),
    .A(\mac1.total_sum[14] ),
    .B(\mac2.total_sum[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5643_ (.A(\mac1.total_sum[14] ),
    .B(\mac2.total_sum[14] ),
    .Y(_2355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5644_ (.B(\mac2.total_sum[14] ),
    .A(\mac1.total_sum[14] ),
    .X(_2356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5645_ (.Y(net23),
    .A(_2353_),
    .B(_2356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5646_ (.B1(_2354_),
    .VDD(VPWR),
    .Y(_2357_),
    .VSS(VGND),
    .A1(_2353_),
    .A2(_2355_));
 sg13g2_xnor2_1 _5647_ (.Y(_2358_),
    .A(\mac1.total_sum[15] ),
    .B(\mac2.total_sum[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5648_ (.Y(net24),
    .A(_2357_),
    .B(_2358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5649_ (.B(\mac2.total_sum[0] ),
    .A(\mac1.total_sum[0] ),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5650_ (.A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ),
    .X(_2359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5651_ (.Y(_2360_),
    .A(\DP_1.I_range.out_data[5] ),
    .B(_2359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5652_ (.Y(_2361_),
    .B(\DP_1.Q_range.out_data[5] ),
    .A_N(\DP_1.Q_range.out_data[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _5653_ (.A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ),
    .Y(_2362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _5654_ (.B(\DP_1.Q_range.out_data[3] ),
    .C(_2362_),
    .Y(_2363_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\DP_1.I_range.out_data[3] ));
 sg13g2_nor4_1 _5655_ (.A(\DP_1.I_range.out_data[6] ),
    .B(\DP_1.I_range.out_data[4] ),
    .C(\DP_1.Q_range.out_data[4] ),
    .D(_2363_),
    .Y(_2364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5656_ (.B1(_2364_),
    .VDD(VPWR),
    .Y(_2365_),
    .VSS(VGND),
    .A1(\DP_1.I_range.out_data[5] ),
    .A2(_2359_));
 sg13g2_a21oi_2 _5657_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2365_),
    .Y(_2366_),
    .A2(_2361_),
    .A1(_2360_));
 sg13g2_xor2_1 _5658_ (.B(\DP_1.Q_range.out_data[3] ),
    .A(\DP_1.I_range.out_data[3] ),
    .X(_2367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5659_ (.A(_2359_),
    .B(_2362_),
    .Y(_2368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5660_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2369_),
    .B(_2362_),
    .A(_2359_));
 sg13g2_nor2_2 _5661_ (.A(_2367_),
    .B(net776),
    .Y(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _5662_ (.Y(_2371_),
    .B(\DP_1.I_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\DP_1.Q_range.out_data[2] ));
 sg13g2_xnor2_1 _5663_ (.Y(_2372_),
    .A(_2367_),
    .B(_2371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5664_ (.B1(net771),
    .VDD(VPWR),
    .Y(_2373_),
    .VSS(VGND),
    .A1(\DP_1.matrix[44] ),
    .A2(_2369_));
 sg13g2_a21oi_1 _5665_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2590_),
    .A2(net773),
    .Y(_2374_),
    .B1(_2373_));
 sg13g2_a21o_1 _5666_ (.A2(net764),
    .A1(net269),
    .B1(_2374_),
    .X(_2375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5667_ (.A0(_2590_),
    .A1(_2375_),
    .S(net756),
    .X(_2376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5668_ (.A0(net983),
    .A1(\DP_1.matrix[41] ),
    .S(net775),
    .X(_2377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5669_ (.Y(_2378_),
    .B1(net771),
    .B2(_2377_),
    .A2(net764),
    .A1(net948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5670_ (.Y(_2379_),
    .A(net326),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5671_ (.A(net987),
    .B(net776),
    .Y(_2380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5672_ (.B1(net772),
    .VDD(VPWR),
    .Y(_2381_),
    .VSS(VGND),
    .A1(net972),
    .A2(net774));
 sg13g2_o21ai_1 _5673_ (.B1(_2379_),
    .VDD(VPWR),
    .Y(_2382_),
    .VSS(VGND),
    .A1(_2380_),
    .A2(_2381_));
 sg13g2_mux2_1 _5674_ (.A0(net977),
    .A1(net993),
    .S(net774),
    .X(_2383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5675_ (.Y(_2384_),
    .B1(net770),
    .B2(_2383_),
    .A2(net763),
    .A1(net959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5676_ (.A(net991),
    .B(net776),
    .Y(_2385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5677_ (.Y(_2386_),
    .A(net957),
    .B(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5678_ (.B1(net770),
    .VDD(VPWR),
    .Y(_2387_),
    .VSS(VGND),
    .A1(net975),
    .A2(net774));
 sg13g2_a22oi_1 _5679_ (.Y(_2388_),
    .B1(_2386_),
    .B2(_2387_),
    .A2(_2385_),
    .A1(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5680_ (.Y(_2389_),
    .B(_2388_),
    .A_N(_2384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5681_ (.Y(_2390_),
    .A(net276),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5682_ (.B1(net770),
    .VDD(VPWR),
    .Y(_2391_),
    .VSS(VGND),
    .A1(net973),
    .A2(net773));
 sg13g2_inv_1 _5683_ (.VDD(VPWR),
    .Y(_2392_),
    .A(_2391_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5684_ (.B1(_2392_),
    .VDD(VPWR),
    .Y(_2393_),
    .VSS(VGND),
    .A1(net989),
    .A2(net776));
 sg13g2_a21o_1 _5685_ (.A2(_2393_),
    .A1(_2390_),
    .B1(_2389_),
    .X(_2394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5686_ (.Y(_2395_),
    .B(_2382_),
    .A_N(_2394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5687_ (.Y(_2396_),
    .A(net951),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5688_ (.A(net985),
    .B(net775),
    .Y(_2397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5689_ (.B1(net772),
    .VDD(VPWR),
    .Y(_2398_),
    .VSS(VGND),
    .A1(net970),
    .A2(net773));
 sg13g2_o21ai_1 _5690_ (.B1(_2396_),
    .VDD(VPWR),
    .Y(_2399_),
    .VSS(VGND),
    .A1(_2397_),
    .A2(_2398_));
 sg13g2_nor2b_1 _5691_ (.A(_2395_),
    .B_N(_2399_),
    .Y(_2400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5692_ (.A(_2378_),
    .B_N(_2400_),
    .Y(_2401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5693_ (.A0(net981),
    .A1(\DP_1.matrix[42] ),
    .S(net775),
    .X(_2402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5694_ (.Y(_2403_),
    .B1(net771),
    .B2(_2402_),
    .A2(net764),
    .A1(net278),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5695_ (.Y(_2404_),
    .B(_2401_),
    .A_N(_2403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5696_ (.A0(net979),
    .A1(net962),
    .S(net776),
    .X(_2405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5697_ (.Y(_2406_),
    .B1(net771),
    .B2(_2405_),
    .A2(net764),
    .A1(net270),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5698_ (.B1(net755),
    .VDD(VPWR),
    .Y(_2407_),
    .VSS(VGND),
    .A1(_2404_),
    .A2(_2406_));
 sg13g2_nor2_1 _5699_ (.A(_2375_),
    .B(_2407_),
    .Y(_2408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5700_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2376_),
    .A2(_2407_),
    .Y(_0160_),
    .B1(_2408_));
 sg13g2_o21ai_1 _5701_ (.B1(net771),
    .VDD(VPWR),
    .Y(_2409_),
    .VSS(VGND),
    .A1(\DP_2.matrix[44] ),
    .A2(net773));
 sg13g2_a21oi_1 _5702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2591_),
    .A2(net773),
    .Y(_2410_),
    .B1(_2409_));
 sg13g2_a21o_1 _5703_ (.A2(net764),
    .A1(net275),
    .B1(_2410_),
    .X(_2411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5704_ (.A0(net927),
    .A1(net911),
    .S(net775),
    .X(_2412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5705_ (.Y(_2413_),
    .B1(net771),
    .B2(_2412_),
    .A2(net764),
    .A1(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5706_ (.Y(_2414_),
    .A(net895),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5707_ (.A(net929),
    .B(net775),
    .Y(_2415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5708_ (.B1(net770),
    .VDD(VPWR),
    .Y(_2416_),
    .VSS(VGND),
    .A1(\DP_2.matrix[39] ),
    .A2(net773));
 sg13g2_o21ai_1 _5709_ (.B1(_2414_),
    .VDD(VPWR),
    .Y(_2417_),
    .VSS(VGND),
    .A1(_2415_),
    .A2(_2416_));
 sg13g2_mux2_1 _5710_ (.A0(net924),
    .A1(net937),
    .S(net774),
    .X(_2418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5711_ (.Y(_2419_),
    .B1(net770),
    .B2(_2418_),
    .A2(net763),
    .A1(net277),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5712_ (.A(net932),
    .B(net776),
    .Y(_2420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5713_ (.Y(_2421_),
    .A(net902),
    .B(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5714_ (.B1(net770),
    .VDD(VPWR),
    .Y(_2422_),
    .VSS(VGND),
    .A1(net918),
    .A2(net774));
 sg13g2_a22oi_1 _5715_ (.Y(_2423_),
    .B1(_2421_),
    .B2(_2422_),
    .A2(_2420_),
    .A1(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5716_ (.Y(_2424_),
    .B(_2423_),
    .A_N(_2419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5717_ (.Y(_2425_),
    .A(net897),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5718_ (.B1(net771),
    .VDD(VPWR),
    .Y(_2426_),
    .VSS(VGND),
    .A1(net916),
    .A2(net773));
 sg13g2_inv_1 _5719_ (.VDD(VPWR),
    .Y(_2427_),
    .A(_2426_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5720_ (.B1(_2427_),
    .VDD(VPWR),
    .Y(_2428_),
    .VSS(VGND),
    .A1(net930),
    .A2(net776));
 sg13g2_a21o_1 _5721_ (.A2(_2428_),
    .A1(_2425_),
    .B1(_2424_),
    .X(_2429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5722_ (.Y(_2430_),
    .B(_2417_),
    .A_N(_2429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5723_ (.Y(_2431_),
    .A(net893),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5724_ (.A(net928),
    .B(net775),
    .Y(_2432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5725_ (.B1(net771),
    .VDD(VPWR),
    .Y(_2433_),
    .VSS(VGND),
    .A1(\DP_2.matrix[40] ),
    .A2(net773));
 sg13g2_o21ai_1 _5726_ (.B1(_2431_),
    .VDD(VPWR),
    .Y(_2434_),
    .VSS(VGND),
    .A1(_2432_),
    .A2(_2433_));
 sg13g2_nor2b_1 _5727_ (.A(_2430_),
    .B_N(_2434_),
    .Y(_2435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5728_ (.A(_2413_),
    .B_N(_2435_),
    .Y(_2436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5729_ (.A0(net926),
    .A1(net909),
    .S(net775),
    .X(_2437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5730_ (.Y(_2438_),
    .B1(net772),
    .B2(_2437_),
    .A2(net764),
    .A1(net280),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5731_ (.Y(_2439_),
    .B(_2436_),
    .A_N(_2438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5732_ (.A0(net925),
    .A1(net907),
    .S(net775),
    .X(_2440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5733_ (.Y(_2441_),
    .B1(net772),
    .B2(_2440_),
    .A2(net764),
    .A1(net888),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5734_ (.A0(_2591_),
    .A1(_2411_),
    .S(net755),
    .X(_2442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5735_ (.B1(net756),
    .VDD(VPWR),
    .Y(_2443_),
    .VSS(VGND),
    .A1(_2439_),
    .A2(_2441_));
 sg13g2_nor2_1 _5736_ (.A(_2411_),
    .B(_2443_),
    .Y(_2444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5737_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2442_),
    .A2(_2443_),
    .Y(_0163_),
    .B1(_2444_));
 sg13g2_nand2b_1 _5738_ (.Y(_2445_),
    .B(\DP_3.I_range.out_data[2] ),
    .A_N(\DP_3.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5739_ (.B(\DP_3.Q_range.out_data[3] ),
    .A(\DP_3.I_range.out_data[3] ),
    .X(_2446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5740_ (.Y(_2447_),
    .A(_2445_),
    .B(_2446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5741_ (.Y(_2448_),
    .A(\DP_3.I_range.out_data[2] ),
    .B(\DP_3.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5742_ (.B(\DP_3.Q_range.out_data[2] ),
    .A(\DP_3.I_range.out_data[2] ),
    .X(_2449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5743_ (.B1(net768),
    .VDD(VPWR),
    .Y(_2450_),
    .VSS(VGND),
    .A1(net1001),
    .A2(net777));
 sg13g2_a21oi_1 _5744_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2592_),
    .A2(net777),
    .Y(_2451_),
    .B1(_2450_));
 sg13g2_nor4_1 _5745_ (.A(\DP_3.Q_range.out_data[2] ),
    .B(_2589_),
    .C(\DP_3.Q_range.out_data[4] ),
    .D(\DP_3.Q_range.out_data[6] ),
    .Y(_2452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5746_ (.A(\DP_3.I_range.out_data[6] ),
    .B(\DP_3.I_range.out_data[2] ),
    .C(_2588_),
    .D(\DP_3.I_range.out_data[4] ),
    .Y(_2453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5747_ (.A(_2446_),
    .B(net778),
    .Y(_2454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5748_ (.Y(_2455_),
    .A(net274),
    .B(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5749_ (.A(net862),
    .B(net779),
    .Y(_2456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5750_ (.B1(net768),
    .VDD(VPWR),
    .Y(_2457_),
    .VSS(VGND),
    .A1(net876),
    .A2(net777));
 sg13g2_o21ai_1 _5751_ (.B1(_2455_),
    .VDD(VPWR),
    .Y(_2458_),
    .VSS(VGND),
    .A1(_2456_),
    .A2(_2457_));
 sg13g2_mux2_1 _5752_ (.A0(net865),
    .A1(net880),
    .S(net780),
    .X(_2459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5753_ (.Y(_2460_),
    .B1(_2459_),
    .B2(net769),
    .A2(net765),
    .A1(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5754_ (.A0(net871),
    .A1(net886),
    .S(net780),
    .X(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5755_ (.Y(_2462_),
    .B1(_2461_),
    .B2(net767),
    .A2(net765),
    .A1(net854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5756_ (.Y(_2463_),
    .A(_2446_),
    .B(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5757_ (.A(net884),
    .B(_2463_),
    .Y(_2464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5758_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net869),
    .A2(net767),
    .Y(_2465_),
    .B1(net780));
 sg13g2_nor2_1 _5759_ (.A(net852),
    .B(net767),
    .Y(_2466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5760_ (.A(_2464_),
    .B(_2465_),
    .C(_2466_),
    .Y(_2467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5761_ (.A(_2462_),
    .B_N(_2467_),
    .Y(_2468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5762_ (.A0(net867),
    .A1(net882),
    .S(net780),
    .X(_2469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5763_ (.Y(_2470_),
    .B1(_2469_),
    .B2(net767),
    .A2(net765),
    .A1(net851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5764_ (.A(_2470_),
    .B_N(_2468_),
    .Y(_2471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5765_ (.Y(_2472_),
    .B(_2471_),
    .A_N(_2460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5766_ (.Y(_2473_),
    .A(net271),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5767_ (.A(net863),
    .B(net779),
    .Y(_2474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5768_ (.B1(net767),
    .VDD(VPWR),
    .Y(_2475_),
    .VSS(VGND),
    .A1(net878),
    .A2(net778));
 sg13g2_o21ai_1 _5769_ (.B1(_2473_),
    .VDD(VPWR),
    .Y(_2476_),
    .VSS(VGND),
    .A1(_2474_),
    .A2(_2475_));
 sg13g2_nand2b_1 _5770_ (.Y(_2477_),
    .B(_2476_),
    .A_N(_2472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5771_ (.Y(_2478_),
    .B(_2458_),
    .A_N(_2477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5772_ (.Y(_2479_),
    .A(net843),
    .B(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5773_ (.A(net860),
    .B(net779),
    .Y(_2480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5774_ (.B1(net769),
    .VDD(VPWR),
    .Y(_2481_),
    .VSS(VGND),
    .A1(net874),
    .A2(net777));
 sg13g2_o21ai_1 _5775_ (.B1(_2479_),
    .VDD(VPWR),
    .Y(_2482_),
    .VSS(VGND),
    .A1(_2480_),
    .A2(_2481_));
 sg13g2_nor2b_1 _5776_ (.A(_2478_),
    .B_N(_2482_),
    .Y(_2483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5777_ (.A0(net857),
    .A1(net873),
    .S(_2448_),
    .X(_2484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5778_ (.Y(_2485_),
    .B1(_2484_),
    .B2(net768),
    .A2(net766),
    .A1(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5779_ (.Y(_2486_),
    .B(_2483_),
    .A_N(_2485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5780_ (.B(\DP_3.Q_range.out_data[3] ),
    .C(_2452_),
    .A(_2587_),
    .Y(_2487_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2453_));
 sg13g2_nor2_1 _5781_ (.A(_2451_),
    .B(net760),
    .Y(_2488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5782_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1001),
    .A2(net760),
    .Y(_2489_),
    .B1(_2488_));
 sg13g2_nand2b_1 _5783_ (.Y(_2490_),
    .B(_2486_),
    .A_N(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5784_ (.A(_2451_),
    .B(_2490_),
    .Y(_2491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2489_),
    .A2(_2490_),
    .Y(_0166_),
    .B1(_2491_));
 sg13g2_o21ai_1 _5786_ (.B1(net768),
    .VDD(VPWR),
    .Y(_2492_),
    .VSS(VGND),
    .A1(net996),
    .A2(net777));
 sg13g2_a21oi_1 _5787_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2593_),
    .A2(net777),
    .Y(_2493_),
    .B1(_2492_));
 sg13g2_nand2_1 _5788_ (.Y(_2494_),
    .A(net786),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5789_ (.A(net806),
    .B(net779),
    .Y(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5790_ (.B1(net768),
    .VDD(VPWR),
    .Y(_2496_),
    .VSS(VGND),
    .A1(net822),
    .A2(net777));
 sg13g2_o21ai_1 _5791_ (.B1(_2494_),
    .VDD(VPWR),
    .Y(_2497_),
    .VSS(VGND),
    .A1(_2495_),
    .A2(_2496_));
 sg13g2_mux2_1 _5792_ (.A0(net809),
    .A1(net825),
    .S(net779),
    .X(_2498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5793_ (.Y(_2499_),
    .B1(_2498_),
    .B2(net769),
    .A2(net765),
    .A1(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5794_ (.A0(net819),
    .A1(net833),
    .S(net780),
    .X(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5795_ (.Y(_2501_),
    .B1(_2500_),
    .B2(net767),
    .A2(net765),
    .A1(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5796_ (.A(net829),
    .B(_2463_),
    .Y(_2502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5797_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net813),
    .A2(net767),
    .Y(_2503_),
    .B1(net780));
 sg13g2_nor2_1 _5798_ (.A(net796),
    .B(net767),
    .Y(_2504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5799_ (.A(_2502_),
    .B(_2503_),
    .C(_2504_),
    .Y(_2505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5800_ (.A(_2501_),
    .B_N(_2505_),
    .Y(_2506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5801_ (.A0(net811),
    .A1(net827),
    .S(net780),
    .X(_2507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5802_ (.Y(_2508_),
    .B1(_2507_),
    .B2(net769),
    .A2(net765),
    .A1(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5803_ (.A(_2508_),
    .B_N(_2506_),
    .Y(_2509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5804_ (.Y(_2510_),
    .B(_2509_),
    .A_N(_2499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5805_ (.Y(_2511_),
    .A(net788),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5806_ (.A(net808),
    .B(net779),
    .Y(_2512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5807_ (.B1(net768),
    .VDD(VPWR),
    .Y(_2513_),
    .VSS(VGND),
    .A1(net824),
    .A2(net777));
 sg13g2_o21ai_1 _5808_ (.B1(_2511_),
    .VDD(VPWR),
    .Y(_2514_),
    .VSS(VGND),
    .A1(_2512_),
    .A2(_2513_));
 sg13g2_nand2b_1 _5809_ (.Y(_2515_),
    .B(_2514_),
    .A_N(_2510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5810_ (.Y(_2516_),
    .B(_2497_),
    .A_N(_2515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5811_ (.Y(_2517_),
    .A(net784),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5812_ (.A(net804),
    .B(net779),
    .Y(_2518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5813_ (.B1(net768),
    .VDD(VPWR),
    .Y(_2519_),
    .VSS(VGND),
    .A1(net821),
    .A2(net778));
 sg13g2_o21ai_1 _5814_ (.B1(_2517_),
    .VDD(VPWR),
    .Y(_2520_),
    .VSS(VGND),
    .A1(_2518_),
    .A2(_2519_));
 sg13g2_nor2b_1 _5815_ (.A(_2516_),
    .B_N(_2520_),
    .Y(_2521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5816_ (.A0(net802),
    .A1(net820),
    .S(net779),
    .X(_2522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5817_ (.Y(_2523_),
    .B1(_2522_),
    .B2(net768),
    .A2(net766),
    .A1(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5818_ (.Y(_2524_),
    .B(_2521_),
    .A_N(_2523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5819_ (.A(net760),
    .B(_2493_),
    .Y(_2525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net996),
    .A2(net760),
    .Y(_2526_),
    .B1(_2525_));
 sg13g2_nand2b_1 _5821_ (.Y(_2527_),
    .B(_2524_),
    .A_N(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5822_ (.A(_2493_),
    .B(_2527_),
    .Y(_2528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2526_),
    .A2(_2527_),
    .Y(_0169_),
    .B1(_2528_));
 sg13g2_xor2_1 _5824_ (.B(net754),
    .A(net993),
    .X(_0172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5825_ (.A(net991),
    .B(net754),
    .Y(_2529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5826_ (.B(_2388_),
    .A(_2384_),
    .X(_2530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5827_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net754),
    .A2(_2530_),
    .Y(_0173_),
    .B1(_2529_));
 sg13g2_nor2_1 _5828_ (.A(net989),
    .B(net753),
    .Y(_2531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5829_ (.B(_2390_),
    .C(_2393_),
    .A(_2389_),
    .Y(_2532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5830_ (.Y(_2533_),
    .A(_2394_),
    .B(_2532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5831_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net754),
    .A2(_2533_),
    .Y(_0174_),
    .B1(_2531_));
 sg13g2_nor2_1 _5832_ (.A(net987),
    .B(net753),
    .Y(_2534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5833_ (.B(_2394_),
    .A(_2382_),
    .X(_2535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5834_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net753),
    .A2(_2535_),
    .Y(_0175_),
    .B1(_2534_));
 sg13g2_nor2_1 _5835_ (.A(net985),
    .B(net753),
    .Y(_2536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5836_ (.B(_2399_),
    .A(_2395_),
    .X(_2537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5837_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net753),
    .A2(_2537_),
    .Y(_0176_),
    .B1(_2536_));
 sg13g2_nor2_1 _5838_ (.A(net983),
    .B(net756),
    .Y(_2538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5839_ (.B(_2400_),
    .A(_2378_),
    .X(_2539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5840_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net756),
    .A2(_2539_),
    .Y(_0177_),
    .B1(_2538_));
 sg13g2_nor2_1 _5841_ (.A(net981),
    .B(net755),
    .Y(_2540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5842_ (.B(_2403_),
    .A(_2401_),
    .X(_2541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5843_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net756),
    .A2(_2541_),
    .Y(_0178_),
    .B1(_2540_));
 sg13g2_nand2b_1 _5844_ (.Y(_2542_),
    .B(net979),
    .A_N(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5845_ (.A(_2404_),
    .B(_2406_),
    .X(_2543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5846_ (.B1(_2542_),
    .VDD(VPWR),
    .Y(_0179_),
    .VSS(VGND),
    .A1(_2407_),
    .A2(_2543_));
 sg13g2_xor2_1 _5847_ (.B(net754),
    .A(net937),
    .X(_0196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5848_ (.A(net932),
    .B(net754),
    .Y(_2544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5849_ (.B(_2423_),
    .A(_2419_),
    .X(_2545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net754),
    .A2(_2545_),
    .Y(_0197_),
    .B1(_2544_));
 sg13g2_nor2_1 _5851_ (.A(net930),
    .B(net753),
    .Y(_2546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5852_ (.B(_2425_),
    .C(_2428_),
    .A(_2424_),
    .Y(_2547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5853_ (.Y(_2548_),
    .A(_2429_),
    .B(_2547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net757),
    .A2(_2548_),
    .Y(_0198_),
    .B1(_2546_));
 sg13g2_nor2_1 _5855_ (.A(net929),
    .B(net753),
    .Y(_2549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5856_ (.B(_2429_),
    .A(_2417_),
    .X(_2550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5857_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net753),
    .A2(_2550_),
    .Y(_0199_),
    .B1(_2549_));
 sg13g2_nor2_1 _5858_ (.A(net928),
    .B(net757),
    .Y(_2551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5859_ (.B(_2434_),
    .A(_2430_),
    .X(_2552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net757),
    .A2(_2552_),
    .Y(_0200_),
    .B1(net432));
 sg13g2_nor2_1 _5861_ (.A(net927),
    .B(net755),
    .Y(_2553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5862_ (.B(_2435_),
    .A(_2413_),
    .X(_2554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5863_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net755),
    .A2(_2554_),
    .Y(_0201_),
    .B1(_2553_));
 sg13g2_nor2_1 _5864_ (.A(net926),
    .B(net755),
    .Y(_2555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5865_ (.B(_2438_),
    .A(_2436_),
    .X(_2556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net755),
    .A2(_2556_),
    .Y(_0202_),
    .B1(_2555_));
 sg13g2_nand2b_1 _5867_ (.Y(_2557_),
    .B(net925),
    .A_N(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5868_ (.A(_2439_),
    .B(_2441_),
    .X(_2558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5869_ (.B1(_2557_),
    .VDD(VPWR),
    .Y(_0203_),
    .VSS(VGND),
    .A1(_2443_),
    .A2(_2558_));
 sg13g2_xnor2_1 _5870_ (.Y(_0220_),
    .A(net886),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5871_ (.B(_2467_),
    .A(_2462_),
    .X(_2559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5872_ (.Y(_2560_),
    .A(net884),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5873_ (.B1(_2560_),
    .VDD(VPWR),
    .Y(_0221_),
    .VSS(VGND),
    .A1(net758),
    .A2(_2559_));
 sg13g2_xor2_1 _5874_ (.B(_2470_),
    .A(_2468_),
    .X(_2561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5875_ (.Y(_2562_),
    .A(net882),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5876_ (.B1(_2562_),
    .VDD(VPWR),
    .Y(_0222_),
    .VSS(VGND),
    .A1(net758),
    .A2(_2561_));
 sg13g2_xor2_1 _5877_ (.B(_2471_),
    .A(_2460_),
    .X(_2563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5878_ (.Y(_2564_),
    .A(net880),
    .B(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5879_ (.B1(_2564_),
    .VDD(VPWR),
    .Y(_0223_),
    .VSS(VGND),
    .A1(net759),
    .A2(_2563_));
 sg13g2_nand2_1 _5880_ (.Y(_2565_),
    .A(net878),
    .B(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5881_ (.B(_2476_),
    .A(_2472_),
    .X(_2566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5882_ (.B1(_2565_),
    .VDD(VPWR),
    .Y(_0224_),
    .VSS(VGND),
    .A1(net759),
    .A2(_2566_));
 sg13g2_nand2_1 _5883_ (.Y(_2567_),
    .A(net876),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5884_ (.B(_2477_),
    .A(_2458_),
    .X(_2568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5885_ (.B1(_2567_),
    .VDD(VPWR),
    .Y(_0225_),
    .VSS(VGND),
    .A1(net761),
    .A2(_2568_));
 sg13g2_xor2_1 _5886_ (.B(_2482_),
    .A(_2478_),
    .X(_2569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5887_ (.Y(_2570_),
    .A(net874),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5888_ (.B1(_2570_),
    .VDD(VPWR),
    .Y(_0226_),
    .VSS(VGND),
    .A1(net761),
    .A2(_2569_));
 sg13g2_nand2_1 _5889_ (.Y(_2571_),
    .A(net873),
    .B(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5890_ (.A(_2483_),
    .B_N(_2485_),
    .Y(_2572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5891_ (.B1(net397),
    .VDD(VPWR),
    .Y(_0227_),
    .VSS(VGND),
    .A1(_2490_),
    .A2(_2572_));
 sg13g2_xnor2_1 _5892_ (.Y(_0244_),
    .A(net833),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5893_ (.B(_2505_),
    .A(_2501_),
    .X(_2573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5894_ (.Y(_2574_),
    .A(net829),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5895_ (.B1(_2574_),
    .VDD(VPWR),
    .Y(_0245_),
    .VSS(VGND),
    .A1(net758),
    .A2(_2573_));
 sg13g2_xor2_1 _5896_ (.B(_2508_),
    .A(_2506_),
    .X(_2575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5897_ (.Y(_2576_),
    .A(net827),
    .B(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5898_ (.B1(_2576_),
    .VDD(VPWR),
    .Y(_0246_),
    .VSS(VGND),
    .A1(net759),
    .A2(_2575_));
 sg13g2_xor2_1 _5899_ (.B(_2509_),
    .A(_2499_),
    .X(_2577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5900_ (.Y(_2578_),
    .A(net825),
    .B(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5901_ (.B1(_2578_),
    .VDD(VPWR),
    .Y(_0247_),
    .VSS(VGND),
    .A1(net762),
    .A2(_2577_));
 sg13g2_nand2_1 _5902_ (.Y(_2579_),
    .A(net824),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5903_ (.B(_2514_),
    .A(_2510_),
    .X(_2580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5904_ (.B1(_2579_),
    .VDD(VPWR),
    .Y(_0248_),
    .VSS(VGND),
    .A1(net761),
    .A2(_2580_));
 sg13g2_nand2_1 _5905_ (.Y(_2581_),
    .A(net822),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5906_ (.B(_2515_),
    .A(_2497_),
    .X(_2582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5907_ (.B1(_2581_),
    .VDD(VPWR),
    .Y(_0249_),
    .VSS(VGND),
    .A1(net761),
    .A2(_2582_));
 sg13g2_xor2_1 _5908_ (.B(_2520_),
    .A(_2516_),
    .X(_2583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5909_ (.Y(_2584_),
    .A(net821),
    .B(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5910_ (.B1(_2584_),
    .VDD(VPWR),
    .Y(_0250_),
    .VSS(VGND),
    .A1(net760),
    .A2(_2583_));
 sg13g2_nand2_1 _5911_ (.Y(_2585_),
    .A(net820),
    .B(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5912_ (.A(_2521_),
    .B_N(_2523_),
    .Y(_2586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5913_ (.B1(_2585_),
    .VDD(VPWR),
    .Y(_0251_),
    .VSS(VGND),
    .A1(_2527_),
    .A2(_2586_));
 sg13g2_buf_1 _5914_ (.A(net1009),
    .X(_0161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5915_ (.A(net269),
    .X(_0162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5916_ (.A(net1004),
    .X(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5917_ (.A(net275),
    .X(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5918_ (.A(net999),
    .X(_0167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5919_ (.A(net997),
    .X(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5920_ (.A(net273),
    .X(_0170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5921_ (.A(net272),
    .X(_0171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5922_ (.A(net281),
    .X(_0180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5923_ (.A(net976),
    .X(_0181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5924_ (.A(net974),
    .X(_0182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5925_ (.A(net971),
    .X(_0183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5926_ (.A(net968),
    .X(_0184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5927_ (.A(net966),
    .X(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5928_ (.A(net963),
    .X(_0186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5929_ (.A(net961),
    .X(_0187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5930_ (.A(net959),
    .X(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5931_ (.A(net957),
    .X(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5932_ (.A(net276),
    .X(_0190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5933_ (.A(net953),
    .X(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5934_ (.A(net951),
    .X(_0192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5935_ (.A(net948),
    .X(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5936_ (.A(net278),
    .X(_0194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5937_ (.A(net270),
    .X(_0195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5938_ (.A(net923),
    .X(_0204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5939_ (.A(net920),
    .X(_0205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5940_ (.A(net916),
    .X(_0206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5941_ (.A(net914),
    .X(_0207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5942_ (.A(net912),
    .X(_0208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5943_ (.A(net910),
    .X(_0209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5944_ (.A(net908),
    .X(_0210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5945_ (.A(net906),
    .X(_0211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5946_ (.A(net277),
    .X(_0212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5947_ (.A(net902),
    .X(_0213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5948_ (.A(net897),
    .X(_0214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5949_ (.A(net895),
    .X(_0215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5950_ (.A(net893),
    .X(_0216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5951_ (.A(net891),
    .X(_0217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5952_ (.A(net280),
    .X(_0218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5953_ (.A(net888),
    .X(_0219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5954_ (.A(net871),
    .X(_0228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5955_ (.A(net869),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5956_ (.A(net867),
    .X(_0230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5957_ (.A(net865),
    .X(_0231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5958_ (.A(net863),
    .X(_0232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5959_ (.A(net861),
    .X(_0233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5960_ (.A(net858),
    .X(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5961_ (.A(net856),
    .X(_0235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5962_ (.A(net279),
    .X(_0236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5963_ (.A(net853),
    .X(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5964_ (.A(net851),
    .X(_0238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5965_ (.A(net849),
    .X(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5966_ (.A(net271),
    .X(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5967_ (.A(net274),
    .X(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5968_ (.A(net843),
    .X(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5969_ (.A(net840),
    .X(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5970_ (.A(net819),
    .X(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5971_ (.A(net813),
    .X(_0253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5972_ (.A(net811),
    .X(_0254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5973_ (.A(net809),
    .X(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5974_ (.A(net808),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5975_ (.A(net805),
    .X(_0257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5976_ (.A(net803),
    .X(_0258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5977_ (.A(net801),
    .X(_0259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5978_ (.A(net800),
    .X(_0260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5979_ (.A(net796),
    .X(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5980_ (.A(net792),
    .X(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5981_ (.A(net790),
    .X(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5982_ (.A(net788),
    .X(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5983_ (.A(net786),
    .X(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5984_ (.A(net784),
    .X(_0266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5985_ (.A(net782),
    .X(_0267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_2 _5986_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net9),
    .Q(\DP_3.Q_range.out_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5987_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net10),
    .Q(\DP_3.Q_range.out_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5988_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net11),
    .Q(\DP_3.Q_range.out_data[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5989_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_3.Q_range.data_plus_4[6] ),
    .Q(\DP_3.Q_range.out_data[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5990_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net12),
    .Q(\DP_3.Q_range.out_data[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5991_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _5992_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _5993_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\mac1.products_ff[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _5994_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(\mac1.products_ff[3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _5995_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\mac1.products_ff[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _5996_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0105_),
    .Q(\mac1.products_ff[5] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _5997_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\mac1.products_ff[6] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _5998_ (.RESET_B(net1069),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0113_),
    .Q(\mac1.products_ff[7] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _5999_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0114_),
    .Q(\mac1.products_ff[8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6000_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\mac1.products_ff[9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6001_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0106_),
    .Q(\mac1.products_ff[10] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6002_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\mac1.products_ff[11] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6003_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0108_),
    .Q(\mac1.products_ff[12] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6004_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\mac1.products_ff[13] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6005_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\mac1.products_ff[14] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6006_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\mac1.products_ff[15] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6007_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\mac1.products_ff[68] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6008_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\mac1.products_ff[69] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6009_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\mac1.products_ff[70] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6010_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\mac1.products_ff[71] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6011_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\mac1.products_ff[72] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6012_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\mac1.products_ff[73] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6013_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\mac1.products_ff[74] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6014_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\mac1.products_ff[75] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6015_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\mac1.products_ff[76] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6016_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\mac1.products_ff[77] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6017_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\mac1.products_ff[78] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6018_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\mac1.products_ff[79] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6019_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0119_),
    .Q(\mac1.products_ff[80] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6020_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\mac1.products_ff[81] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6021_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\mac1.products_ff[82] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6022_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\mac1.products_ff[83] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6023_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net446),
    .Q(\DP_1.matrix[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6024_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\DP_1.matrix[44] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6025_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\DP_1.matrix[80] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6026_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\DP_2.matrix[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6027_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\DP_2.matrix[44] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6028_ (.RESET_B(net1048),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\DP_2.matrix[80] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6029_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\DP_3.matrix[8] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6030_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\DP_3.matrix[44] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6031_ (.RESET_B(net1037),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\DP_3.matrix[80] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6032_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0169_),
    .Q(\DP_4.matrix[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6033_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\DP_4.matrix[44] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6034_ (.RESET_B(net1037),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\DP_4.matrix[80] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6035_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6036_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6037_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\DP_1.matrix[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6038_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\DP_1.matrix[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6039_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\DP_1.matrix[4] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6040_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\DP_1.matrix[5] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6041_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\DP_1.matrix[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6042_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\DP_1.matrix[7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6043_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\DP_1.matrix[36] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6044_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0181_),
    .Q(\DP_1.matrix[37] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6045_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0182_),
    .Q(\DP_1.matrix[38] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6046_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0183_),
    .Q(\DP_1.matrix[39] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6047_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\DP_1.matrix[40] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6048_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0185_),
    .Q(\DP_1.matrix[41] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6049_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\mac1.products_ff[136] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6050_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\DP_1.matrix[42] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6051_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(\DP_1.matrix[43] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6052_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\mac1.products_ff[137] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6053_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0188_),
    .Q(\DP_1.matrix[72] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6054_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0189_),
    .Q(\DP_1.matrix[73] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6055_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\mac1.products_ff[138] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6056_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\DP_1.matrix[74] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6057_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\DP_1.matrix[75] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6058_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0067_),
    .Q(\mac1.products_ff[139] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6059_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\DP_1.matrix[76] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6060_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\DP_1.matrix[77] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6061_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\mac1.products_ff[140] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _6062_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\DP_1.matrix[78] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6063_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0195_),
    .Q(\DP_1.matrix[79] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6064_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\mac1.products_ff[141] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6065_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0196_),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6066_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0197_),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6067_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\mac1.products_ff[142] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6068_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net389),
    .Q(\DP_2.matrix[2] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6069_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0199_),
    .Q(\DP_2.matrix[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6070_ (.RESET_B(net1015),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\mac1.products_ff[143] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6071_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0200_),
    .Q(\DP_2.matrix[4] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6072_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0201_),
    .Q(\DP_2.matrix[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6073_ (.RESET_B(net1015),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0103_),
    .Q(\mac1.products_ff[144] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6074_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0202_),
    .Q(\DP_2.matrix[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6075_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0203_),
    .Q(\DP_2.matrix[7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6076_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\mac1.products_ff[145] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6077_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0204_),
    .Q(\DP_2.matrix[36] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6078_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0205_),
    .Q(\DP_2.matrix[37] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6079_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\mac1.products_ff[146] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6080_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0206_),
    .Q(\DP_2.matrix[38] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6081_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\DP_2.matrix[39] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6082_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\mac1.products_ff[147] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6083_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0208_),
    .Q(\DP_2.matrix[40] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6084_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0209_),
    .Q(\DP_2.matrix[41] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6085_ (.RESET_B(net1021),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0097_),
    .Q(\mac1.products_ff[148] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6086_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0210_),
    .Q(\DP_2.matrix[42] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6087_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0211_),
    .Q(\DP_2.matrix[43] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6088_ (.RESET_B(net1025),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\mac1.products_ff[149] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6089_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0212_),
    .Q(\DP_2.matrix[72] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6090_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0213_),
    .Q(\DP_2.matrix[73] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6091_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\mac1.products_ff[150] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6092_ (.RESET_B(net1063),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0214_),
    .Q(\DP_2.matrix[74] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6093_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0215_),
    .Q(\DP_2.matrix[75] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6094_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\mac1.products_ff[151] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6095_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0216_),
    .Q(\DP_2.matrix[76] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6096_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0217_),
    .Q(\DP_2.matrix[77] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6097_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net89),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6098_ (.RESET_B(net1048),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0218_),
    .Q(\DP_2.matrix[78] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6099_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0219_),
    .Q(\DP_2.matrix[79] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6100_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net198),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6101_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0220_),
    .Q(\DP_3.matrix[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6102_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0221_),
    .Q(\DP_3.matrix[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6103_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net57),
    .Q(\mac1.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6104_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\DP_3.matrix[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6105_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\DP_3.matrix[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6106_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net68),
    .Q(\mac1.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6107_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0224_),
    .Q(\DP_3.matrix[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6108_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0225_),
    .Q(\DP_3.matrix[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6109_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net204),
    .Q(\mac1.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _6110_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\DP_3.matrix[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6111_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\DP_3.matrix[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6112_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net64),
    .Q(\mac1.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6113_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0228_),
    .Q(\DP_3.matrix[36] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6114_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0229_),
    .Q(\DP_3.matrix[37] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6115_ (.RESET_B(net1069),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net147),
    .Q(\mac1.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6116_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0230_),
    .Q(\DP_3.matrix[38] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6117_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0231_),
    .Q(\DP_3.matrix[39] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6118_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net230),
    .Q(\mac1.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6119_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0232_),
    .Q(\DP_3.matrix[40] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6120_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0233_),
    .Q(\DP_3.matrix[41] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6121_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net61),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6122_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0234_),
    .Q(\DP_3.matrix[42] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6123_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0235_),
    .Q(\DP_3.matrix[43] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6124_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net65),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6125_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0236_),
    .Q(\DP_3.matrix[72] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6126_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0237_),
    .Q(\DP_3.matrix[73] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6127_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net98),
    .Q(\mac1.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6128_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0238_),
    .Q(\DP_3.matrix[74] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6129_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0239_),
    .Q(\DP_3.matrix[75] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6130_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net99),
    .Q(\mac1.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6131_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0240_),
    .Q(\DP_3.matrix[76] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6132_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\DP_3.matrix[77] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6133_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net150),
    .Q(\mac1.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6134_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0242_),
    .Q(\DP_3.matrix[78] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6135_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0243_),
    .Q(\DP_3.matrix[79] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6136_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net179),
    .Q(\mac1.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6137_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0244_),
    .Q(\DP_4.matrix[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6138_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\DP_4.matrix[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6139_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net76),
    .Q(\mac1.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6140_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0246_),
    .Q(\DP_4.matrix[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6141_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net351),
    .Q(\DP_4.matrix[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6142_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net80),
    .Q(\mac1.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6143_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0248_),
    .Q(\DP_4.matrix[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6144_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0249_),
    .Q(\DP_4.matrix[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6145_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0250_),
    .Q(\DP_4.matrix[6] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6146_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0251_),
    .Q(\DP_4.matrix[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6147_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0252_),
    .Q(\DP_4.matrix[36] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6148_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0253_),
    .Q(\DP_4.matrix[37] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6149_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0254_),
    .Q(\DP_4.matrix[38] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6150_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0255_),
    .Q(\DP_4.matrix[39] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6151_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\DP_4.matrix[40] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6152_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0257_),
    .Q(\DP_4.matrix[41] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6153_ (.RESET_B(net1095),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0258_),
    .Q(\DP_4.matrix[42] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6154_ (.RESET_B(net1095),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0259_),
    .Q(\DP_4.matrix[43] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6155_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0260_),
    .Q(\DP_4.matrix[72] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6156_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0261_),
    .Q(\DP_4.matrix[73] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6157_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0262_),
    .Q(\DP_4.matrix[74] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6158_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\DP_4.matrix[75] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6159_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\DP_4.matrix[76] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6160_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0265_),
    .Q(\DP_4.matrix[77] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6161_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0266_),
    .Q(\DP_4.matrix[78] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6162_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0267_),
    .Q(\DP_4.matrix[79] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6163_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net224),
    .Q(\mac1.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6164_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net92),
    .Q(\mac1.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6165_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net231),
    .Q(\mac1.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6166_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net134),
    .Q(\mac1.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6167_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net86),
    .Q(\mac1.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6168_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net177),
    .Q(\mac1.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6169_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net237),
    .Q(\mac1.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6170_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net152),
    .Q(\mac1.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6171_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net240),
    .Q(\mac1.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6172_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net149),
    .Q(\mac1.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6173_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net247),
    .Q(\mac1.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6174_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net257),
    .Q(\mac1.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6175_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net232),
    .Q(\mac1.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6176_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net210),
    .Q(\mac1.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6177_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net75),
    .Q(\mac1.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6178_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net60),
    .Q(\mac1.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6179_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net146),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6180_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net205),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6181_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net114),
    .Q(\mac1.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6182_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net187),
    .Q(\mac1.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6183_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net101),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6184_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net157),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6185_ (.RESET_B(net1069),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net162),
    .Q(\mac1.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6186_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net127),
    .Q(\mac1.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6187_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net151),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6188_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net71),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6189_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net135),
    .Q(\mac1.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6190_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net49),
    .Q(\mac1.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6191_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net94),
    .Q(\mac1.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6192_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net110),
    .Q(\mac1.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6193_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net103),
    .Q(\mac1.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6194_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net100),
    .Q(\mac1.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6195_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net197),
    .Q(\mac1.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6196_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net96),
    .Q(\mac1.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6197_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net131),
    .Q(\mac1.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6198_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net116),
    .Q(\mac1.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6199_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net160),
    .Q(\mac1.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _6200_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net41),
    .Q(\mac1.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6201_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net183),
    .Q(\mac1.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6202_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net173),
    .Q(\mac1.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6203_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net192),
    .Q(\mac1.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6204_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net239),
    .Q(\mac1.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6205_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net46),
    .Q(\mac1.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6206_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net221),
    .Q(\mac1.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6207_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net220),
    .Q(\mac1.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6208_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net242),
    .Q(\mac1.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6209_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net217),
    .Q(\mac1.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6210_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net215),
    .Q(\mac1.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6211_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net148),
    .Q(\mac1.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6212_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net126),
    .Q(\mac1.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6213_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net115),
    .Q(\mac1.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6214_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net87),
    .Q(\mac1.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6215_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net172),
    .Q(\mac1.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6216_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net153),
    .Q(\mac1.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6217_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net201),
    .Q(\mac1.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6218_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net193),
    .Q(\mac1.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6219_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net216),
    .Q(\mac1.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6220_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net180),
    .Q(\mac1.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6221_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net207),
    .Q(\mac1.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6222_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net164),
    .Q(\mac1.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6223_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net236),
    .Q(\mac1.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6224_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net170),
    .Q(\mac1.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6225_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net81),
    .Q(\mac1.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6226_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net213),
    .Q(\mac1.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6227_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net196),
    .Q(\mac2.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6228_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net235),
    .Q(\mac2.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6229_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net182),
    .Q(\mac2.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6230_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net84),
    .Q(\mac2.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6231_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net95),
    .Q(\mac2.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6232_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net194),
    .Q(\mac2.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6233_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net190),
    .Q(\mac2.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6234_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net222),
    .Q(\mac2.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6235_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net104),
    .Q(\mac2.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6236_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net42),
    .Q(\mac2.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6237_ (.RESET_B(net1030),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net52),
    .Q(\mac2.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6238_ (.RESET_B(net1029),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net154),
    .Q(\mac2.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6239_ (.RESET_B(net1038),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net128),
    .Q(\mac2.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6240_ (.RESET_B(net1034),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net243),
    .Q(\mac2.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6241_ (.RESET_B(net1032),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net91),
    .Q(\mac2.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6242_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net250),
    .Q(\mac2.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6243_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net136),
    .Q(\mac1.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6244_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net51),
    .Q(\mac1.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6245_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net249),
    .Q(\mac1.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6246_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net161),
    .Q(\mac1.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6247_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net212),
    .Q(\mac1.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6248_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net175),
    .Q(\mac1.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6249_ (.RESET_B(net1014),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net144),
    .Q(\mac1.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6250_ (.RESET_B(net1015),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net166),
    .Q(\mac1.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6251_ (.RESET_B(net1015),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net43),
    .Q(\mac1.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6252_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net259),
    .Q(\mac1.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6253_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net225),
    .Q(\mac1.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6254_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net176),
    .Q(\mac1.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6255_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net202),
    .Q(\mac1.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6256_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net44),
    .Q(\mac1.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6257_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net206),
    .Q(\mac1.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6258_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net102),
    .Q(\mac1.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6259_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net77),
    .Q(\mac2.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6260_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net66),
    .Q(\mac2.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6261_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net252),
    .Q(\mac2.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6262_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net234),
    .Q(\mac2.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6263_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net255),
    .Q(\mac2.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6264_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net185),
    .Q(\mac2.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6265_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net245),
    .Q(\mac2.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6266_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net208),
    .Q(\mac2.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6267_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net132),
    .Q(\mac2.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6268_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net54),
    .Q(\mac2.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6269_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net211),
    .Q(\mac2.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6270_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net209),
    .Q(\mac2.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6271_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net97),
    .Q(\mac2.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6272_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net219),
    .Q(\mac2.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6273_ (.RESET_B(net1032),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net258),
    .Q(\mac2.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6274_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net199),
    .Q(\mac2.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6275_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net181),
    .Q(\mac1.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6276_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net70),
    .Q(\mac1.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6277_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net171),
    .Q(\mac1.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6278_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net260),
    .Q(\mac1.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6279_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net142),
    .Q(\mac1.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6280_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net120),
    .Q(\mac1.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6281_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net106),
    .Q(\mac1.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6282_ (.RESET_B(net1022),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net143),
    .Q(\mac1.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6283_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net74),
    .Q(\mac1.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6284_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net58),
    .Q(\mac1.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6285_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net123),
    .Q(\mac1.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6286_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net53),
    .Q(\mac1.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6287_ (.RESET_B(net1025),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net55),
    .Q(\mac1.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6288_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net158),
    .Q(\mac1.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6289_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net226),
    .Q(\mac1.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6290_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net129),
    .Q(\mac1.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6291_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net266),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6292_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net334),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6293_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net417),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6294_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net496),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6295_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0010_),
    .Q(\mac1.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6296_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0011_),
    .Q(\mac1.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6297_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0012_),
    .Q(\mac1.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6298_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0013_),
    .Q(\mac1.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6299_ (.RESET_B(net1023),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net501),
    .Q(\mac1.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6300_ (.RESET_B(net1019),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0015_),
    .Q(\mac1.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6301_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\mac1.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6302_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\mac1.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6303_ (.RESET_B(net1024),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\mac1.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6304_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net481),
    .Q(\mac1.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6305_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net470),
    .Q(\mac1.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6306_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net287),
    .Q(\mac1.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6307_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net256),
    .Q(\mac2.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6308_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net145),
    .Q(\mac2.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6309_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net169),
    .Q(\mac2.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6310_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net83),
    .Q(\mac2.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6311_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net233),
    .Q(\mac2.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6312_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net251),
    .Q(\mac2.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6313_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net117),
    .Q(\mac2.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6314_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net67),
    .Q(\mac2.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6315_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net137),
    .Q(\mac2.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6316_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net113),
    .Q(\mac2.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6317_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net85),
    .Q(\mac2.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6318_ (.RESET_B(net1029),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net56),
    .Q(\mac2.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6319_ (.RESET_B(net1029),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net82),
    .Q(\mac2.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6320_ (.RESET_B(net1034),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net48),
    .Q(\mac2.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6321_ (.RESET_B(net1034),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net241),
    .Q(\mac2.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6322_ (.RESET_B(net1034),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net174),
    .Q(\mac2.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6323_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net284),
    .Q(\mac1.total_sum[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6324_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net430),
    .Q(\mac1.total_sum[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6325_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net435),
    .Q(\mac1.total_sum[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6326_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net385),
    .Q(\mac1.total_sum[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6327_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net355),
    .Q(\mac1.total_sum[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6328_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net319),
    .Q(\mac1.total_sum[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6329_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net486),
    .Q(\mac1.total_sum[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6330_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net521),
    .Q(\mac1.total_sum[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6331_ (.RESET_B(net1016),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net408),
    .Q(\mac1.total_sum[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6332_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net295),
    .Q(\mac1.total_sum[9] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6333_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net379),
    .Q(\mac1.total_sum[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6334_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net395),
    .Q(\mac1.total_sum[11] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6335_ (.RESET_B(net1018),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net325),
    .Q(\mac1.total_sum[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6336_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net343),
    .Q(\mac1.total_sum[13] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6337_ (.RESET_B(net1018),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net375),
    .Q(\mac1.total_sum[14] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6338_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net411),
    .Q(\mac1.total_sum[15] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6339_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\mac2.products_ff[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6340_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\mac2.products_ff[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6341_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\mac2.products_ff[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6342_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\mac2.products_ff[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6343_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\mac2.products_ff[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6344_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\mac2.products_ff[5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6345_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\mac2.products_ff[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6346_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\mac2.products_ff[7] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6347_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\mac2.products_ff[8] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6348_ (.RESET_B(net1091),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\mac2.products_ff[9] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6349_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\mac2.products_ff[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6350_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\mac2.products_ff[11] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6351_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\mac2.products_ff[12] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6352_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0142_),
    .Q(\mac2.products_ff[13] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6353_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\mac2.products_ff[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6354_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\mac2.products_ff[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6355_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\mac2.products_ff[68] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6356_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\mac2.products_ff[69] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6357_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\mac2.products_ff[70] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6358_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\mac2.products_ff[71] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6359_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\mac2.products_ff[72] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6360_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\mac2.products_ff[73] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6361_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\mac2.products_ff[74] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6362_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\mac2.products_ff[75] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6363_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\mac2.products_ff[76] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6364_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\mac2.products_ff[77] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6365_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\mac2.products_ff[78] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6366_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\mac2.products_ff[79] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6367_ (.RESET_B(net1091),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\mac2.products_ff[80] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6368_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\mac2.products_ff[81] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6369_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\mac2.products_ff[82] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6370_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\mac2.products_ff[83] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6371_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0089_),
    .Q(\mac2.products_ff[136] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6372_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net290),
    .Q(\mac2.products_ff[137] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6373_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\mac2.products_ff[138] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6374_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\mac2.products_ff[139] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6375_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\mac2.products_ff[140] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6376_ (.RESET_B(net1036),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\mac2.products_ff[141] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6377_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\mac2.products_ff[142] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6378_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0157_),
    .Q(\mac2.products_ff[143] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6379_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\mac2.products_ff[144] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6380_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0159_),
    .Q(\mac2.products_ff[145] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6381_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\mac2.products_ff[146] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6382_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\mac2.products_ff[147] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6383_ (.RESET_B(net1033),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\mac2.products_ff[148] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6384_ (.RESET_B(net1032),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\mac2.products_ff[149] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6385_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\mac2.products_ff[150] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6386_ (.RESET_B(net1032),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\mac2.products_ff[151] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6387_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net253),
    .Q(\mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6388_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net45),
    .Q(\mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6389_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net223),
    .Q(\mac2.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6390_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net78),
    .Q(\mac2.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6391_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net195),
    .Q(\mac2.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6392_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net122),
    .Q(\mac2.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6393_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net254),
    .Q(\mac2.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6394_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net248),
    .Q(\mac2.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6395_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net111),
    .Q(\mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6396_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net228),
    .Q(\mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6397_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net184),
    .Q(\mac2.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6398_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net93),
    .Q(\mac2.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6399_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net263),
    .Q(\mac2.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6400_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net261),
    .Q(\mac2.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6401_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net262),
    .Q(\mac2.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6402_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net264),
    .Q(\mac2.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6403_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net163),
    .Q(\mac2.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6404_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net138),
    .Q(\mac2.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6405_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net203),
    .Q(\mac2.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6406_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net79),
    .Q(\mac2.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6407_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net214),
    .Q(\mac2.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6408_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net229),
    .Q(\mac2.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6409_ (.RESET_B(net1071),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net218),
    .Q(\mac2.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6410_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net189),
    .Q(\mac2.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6411_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net186),
    .Q(\mac2.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6412_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net62),
    .Q(\mac2.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6413_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net191),
    .Q(\mac2.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6414_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net112),
    .Q(\mac2.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6415_ (.RESET_B(net1091),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net167),
    .Q(\mac2.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6416_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net165),
    .Q(\mac2.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6417_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net121),
    .Q(\mac2.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6418_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net168),
    .Q(\mac2.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6419_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1),
    .Q(\DP_1.I_range.out_data[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6420_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2),
    .Q(\DP_1.I_range.out_data[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6421_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3),
    .Q(\DP_1.I_range.out_data[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6422_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_1.I_range.data_plus_4[6] ),
    .Q(\DP_1.I_range.out_data[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6423_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net4),
    .Q(\DP_1.I_range.out_data[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6424_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net47),
    .Q(\mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6425_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net244),
    .Q(\mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6426_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net133),
    .Q(\mac2.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6427_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net109),
    .Q(\mac2.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6428_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net90),
    .Q(\mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6429_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net140),
    .Q(\mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6430_ (.RESET_B(net1071),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net108),
    .Q(\mac2.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6431_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net105),
    .Q(\mac2.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6432_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net227),
    .Q(\mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6433_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net200),
    .Q(\mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6434_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net50),
    .Q(\mac2.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6435_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net107),
    .Q(\mac2.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6436_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net238),
    .Q(\mac2.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6437_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net159),
    .Q(\mac2.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6438_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net178),
    .Q(\mac2.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6439_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net124),
    .Q(\mac2.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6440_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net139),
    .Q(\mac2.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6441_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net119),
    .Q(\mac2.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6442_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net155),
    .Q(\mac2.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6443_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net188),
    .Q(\mac2.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6444_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net69),
    .Q(\mac2.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6445_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net72),
    .Q(\mac2.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6446_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net246),
    .Q(\mac2.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6447_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net156),
    .Q(\mac2.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6448_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net88),
    .Q(\mac2.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6449_ (.RESET_B(net1090),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net125),
    .Q(\mac2.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6450_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net73),
    .Q(\mac2.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6451_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net59),
    .Q(\mac2.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6452_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net141),
    .Q(\mac2.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6453_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net130),
    .Q(\mac2.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6454_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net118),
    .Q(\mac2.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6455_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net63),
    .Q(\mac2.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6456_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net268),
    .Q(\mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6457_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net292),
    .Q(\mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6458_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net322),
    .Q(\mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6459_ (.RESET_B(net1062),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net362),
    .Q(\mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6460_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net463),
    .Q(\mac2.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6461_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net450),
    .Q(\mac2.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6462_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net527),
    .Q(\mac2.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6463_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\mac2.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6464_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net508),
    .Q(\mac2.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6465_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\mac2.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6466_ (.RESET_B(net1035),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\mac2.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6467_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\mac2.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6468_ (.RESET_B(net1029),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\mac2.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6469_ (.RESET_B(net1028),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net513),
    .Q(\mac2.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6470_ (.RESET_B(net1034),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\mac2.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6471_ (.RESET_B(net1037),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\mac2.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6472_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net306),
    .Q(\mac2.total_sum[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6473_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net475),
    .Q(\mac2.total_sum[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6474_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net453),
    .Q(\mac2.total_sum[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6475_ (.RESET_B(net1012),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net489),
    .Q(\mac2.total_sum[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6476_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net456),
    .Q(\mac2.total_sum[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6477_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net420),
    .Q(\mac2.total_sum[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6478_ (.RESET_B(net1016),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net460),
    .Q(\mac2.total_sum[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6479_ (.RESET_B(net1013),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net541),
    .Q(\mac2.total_sum[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6480_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net439),
    .Q(\mac2.total_sum[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6481_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net340),
    .Q(\mac2.total_sum[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6482_ (.RESET_B(net1017),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net382),
    .Q(\mac2.total_sum[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6483_ (.RESET_B(net1018),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net426),
    .Q(\mac2.total_sum[11] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6484_ (.RESET_B(net1018),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net313),
    .Q(\mac2.total_sum[12] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6485_ (.RESET_B(net1018),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net401),
    .Q(\mac2.total_sum[13] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6486_ (.RESET_B(net1018),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net349),
    .Q(\mac2.total_sum[14] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6487_ (.RESET_B(net1020),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net369),
    .Q(\mac2.total_sum[15] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6488_ (.RESET_B(net1027),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net5),
    .Q(\DP_1.Q_range.out_data[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6489_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net6),
    .Q(\DP_1.Q_range.out_data[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6490_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net7),
    .Q(\DP_1.Q_range.out_data[4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6491_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_1.Q_range.data_plus_4[6] ),
    .Q(\DP_1.Q_range.out_data[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6492_ (.RESET_B(net1026),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net8),
    .Q(\DP_1.Q_range.out_data[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6493_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net13),
    .Q(\DP_3.I_range.out_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6494_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net14),
    .Q(\DP_3.I_range.out_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6495_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net15),
    .Q(\DP_3.I_range.out_data[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6496_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_3.I_range.data_plus_4[6] ),
    .Q(\DP_3.I_range.out_data[5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6497_ (.RESET_B(net1031),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net16),
    .Q(\DP_3.I_range.out_data[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_tiehi heichips25_SDR_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi heichips25_SDR_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi heichips25_SDR_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi heichips25_SDR_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi heichips25_SDR_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi heichips25_SDR_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi heichips25_SDR_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout754 (.A(net757),
    .X(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout755 (.A(net756),
    .X(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout756 (.A(net757),
    .X(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout757 (.A(_2366_),
    .X(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout758 (.A(net759),
    .X(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout759 (.A(net762),
    .X(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout760 (.A(net762),
    .X(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout761 (.A(net762),
    .X(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout762 (.A(_2487_),
    .X(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout763 (.A(_2370_),
    .X(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout764 (.A(_2370_),
    .X(net764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout765 (.A(net766),
    .X(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout766 (.A(_2454_),
    .X(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout767 (.A(net769),
    .X(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout769 (.A(_2447_),
    .X(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout770 (.A(net772),
    .X(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout771 (.A(net772),
    .X(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout772 (.A(_2372_),
    .X(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout773 (.A(net774),
    .X(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout774 (.A(_2369_),
    .X(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout775 (.A(net776),
    .X(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout776 (.A(_2368_),
    .X(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout777 (.A(net778),
    .X(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout778 (.A(_2449_),
    .X(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout779 (.A(_2448_),
    .X(net779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout780 (.A(_2448_),
    .X(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout781 (.A(net782),
    .X(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout782 (.A(net309),
    .X(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout784 (.A(net315),
    .X(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout785 (.A(net786),
    .X(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout786 (.A(net356),
    .X(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout787 (.A(net788),
    .X(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout788 (.A(net296),
    .X(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout789 (.A(net790),
    .X(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout790 (.A(net300),
    .X(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout792 (.A(net303),
    .X(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout793 (.A(net795),
    .X(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout794 (.A(net796),
    .X(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout795 (.A(net796),
    .X(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout796 (.A(net288),
    .X(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout797 (.A(net798),
    .X(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout798 (.A(net800),
    .X(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout800 (.A(net282),
    .X(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout801 (.A(net802),
    .X(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout802 (.A(net465),
    .X(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout803 (.A(net804),
    .X(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout804 (.A(net467),
    .X(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout806 (.A(net482),
    .X(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout807 (.A(net808),
    .X(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout808 (.A(net314),
    .X(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout809 (.A(net328),
    .X(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout810 (.A(\DP_4.matrix[39] ),
    .X(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout811 (.A(net331),
    .X(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout812 (.A(\DP_4.matrix[38] ),
    .X(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout813 (.A(net330),
    .X(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout814 (.A(net816),
    .X(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout815 (.A(net816),
    .X(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout816 (.A(\DP_4.matrix[37] ),
    .X(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout817 (.A(net818),
    .X(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout818 (.A(\DP_4.matrix[36] ),
    .X(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout819 (.A(net337),
    .X(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout820 (.A(net428),
    .X(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout821 (.A(net413),
    .X(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout822 (.A(net404),
    .X(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout823 (.A(net824),
    .X(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout824 (.A(net344),
    .X(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout825 (.A(net350),
    .X(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout826 (.A(\DP_4.matrix[3] ),
    .X(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout827 (.A(net366),
    .X(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout828 (.A(\DP_4.matrix[2] ),
    .X(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout829 (.A(net359),
    .X(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout830 (.A(\DP_4.matrix[1] ),
    .X(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout832 (.A(\DP_4.matrix[1] ),
    .X(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout833 (.A(net837),
    .X(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout834 (.A(net837),
    .X(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout835 (.A(net837),
    .X(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout836 (.A(net837),
    .X(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout837 (.A(net376),
    .X(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout838 (.A(net840),
    .X(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout839 (.A(net840),
    .X(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout840 (.A(net298),
    .X(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout841 (.A(net843),
    .X(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout842 (.A(net843),
    .X(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout843 (.A(net308),
    .X(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout844 (.A(net845),
    .X(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout845 (.A(\DP_3.matrix[77] ),
    .X(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout846 (.A(net847),
    .X(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout847 (.A(\DP_3.matrix[76] ),
    .X(net847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout848 (.A(\DP_3.matrix[75] ),
    .X(net848),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout849 (.A(net421),
    .X(net849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout850 (.A(net851),
    .X(net850),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout851 (.A(net302),
    .X(net851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout852 (.A(\DP_3.matrix[73] ),
    .X(net852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout853 (.A(net372),
    .X(net853),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout854 (.A(\DP_3.matrix[72] ),
    .X(net854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout855 (.A(net857),
    .X(net855),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout856 (.A(net857),
    .X(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout857 (.A(net447),
    .X(net857),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout858 (.A(net860),
    .X(net858),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout859 (.A(net860),
    .X(net859),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout860 (.A(net472),
    .X(net860),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout861 (.A(net862),
    .X(net861),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout862 (.A(net497),
    .X(net862),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout863 (.A(net864),
    .X(net863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout864 (.A(net492),
    .X(net864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout865 (.A(net866),
    .X(net865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout866 (.A(net473),
    .X(net866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout867 (.A(net327),
    .X(net867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout868 (.A(\DP_3.matrix[38] ),
    .X(net868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout869 (.A(net329),
    .X(net869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout870 (.A(\DP_3.matrix[37] ),
    .X(net870),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout871 (.A(net363),
    .X(net871),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout872 (.A(\DP_3.matrix[7] ),
    .X(net872),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout873 (.A(net396),
    .X(net873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout874 (.A(net386),
    .X(net874),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout875 (.A(\DP_3.matrix[6] ),
    .X(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout876 (.A(net364),
    .X(net876),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout877 (.A(\DP_3.matrix[5] ),
    .X(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout878 (.A(net879),
    .X(net878),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout879 (.A(net517),
    .X(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout880 (.A(net881),
    .X(net880),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout881 (.A(net493),
    .X(net881),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout882 (.A(net883),
    .X(net882),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout883 (.A(net498),
    .X(net883),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout884 (.A(net370),
    .X(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout885 (.A(\DP_3.matrix[1] ),
    .X(net885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout886 (.A(net365),
    .X(net886),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout887 (.A(net888),
    .X(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout888 (.A(net346),
    .X(net888),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout889 (.A(\DP_2.matrix[78] ),
    .X(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout890 (.A(net891),
    .X(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout891 (.A(net357),
    .X(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout892 (.A(net893),
    .X(net892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout893 (.A(net307),
    .X(net893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout894 (.A(net895),
    .X(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout895 (.A(net301),
    .X(net895),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout896 (.A(net897),
    .X(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout897 (.A(net310),
    .X(net897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout898 (.A(net902),
    .X(net898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout899 (.A(net902),
    .X(net899),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout900 (.A(net901),
    .X(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout901 (.A(net902),
    .X(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout902 (.A(net345),
    .X(net902),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout905 (.A(\DP_2.matrix[72] ),
    .X(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout906 (.A(net907),
    .X(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout907 (.A(net464),
    .X(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout908 (.A(net909),
    .X(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout909 (.A(net466),
    .X(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout910 (.A(net911),
    .X(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout911 (.A(net471),
    .X(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout912 (.A(net913),
    .X(net912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout913 (.A(net523),
    .X(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout914 (.A(net915),
    .X(net914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout915 (.A(net504),
    .X(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout916 (.A(net335),
    .X(net916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout917 (.A(\DP_2.matrix[38] ),
    .X(net917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout918 (.A(net442),
    .X(net918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout920 (.A(net921),
    .X(net920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout921 (.A(\DP_2.matrix[37] ),
    .X(net921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout922 (.A(net923),
    .X(net922),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout923 (.A(net391),
    .X(net923),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout924 (.A(net391),
    .X(net924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout925 (.A(net387),
    .X(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout926 (.A(net414),
    .X(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout927 (.A(net422),
    .X(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout928 (.A(net431),
    .X(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout929 (.A(net444),
    .X(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout930 (.A(net388),
    .X(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout931 (.A(\DP_2.matrix[2] ),
    .X(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout932 (.A(net936),
    .X(net932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout934 (.A(net935),
    .X(net934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout935 (.A(net936),
    .X(net935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout936 (.A(net443),
    .X(net936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout937 (.A(net940),
    .X(net937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout940 (.A(net427),
    .X(net940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout941 (.A(net942),
    .X(net941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout942 (.A(net943),
    .X(net942),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout943 (.A(\DP_1.matrix[79] ),
    .X(net943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout944 (.A(net945),
    .X(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout945 (.A(\DP_1.matrix[78] ),
    .X(net945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout946 (.A(net947),
    .X(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout947 (.A(net948),
    .X(net947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout948 (.A(net336),
    .X(net948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout949 (.A(net951),
    .X(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout950 (.A(net951),
    .X(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout951 (.A(net297),
    .X(net951),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout952 (.A(net953),
    .X(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout953 (.A(net326),
    .X(net953),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout954 (.A(net955),
    .X(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout955 (.A(\DP_1.matrix[74] ),
    .X(net955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout956 (.A(net957),
    .X(net956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout957 (.A(net304),
    .X(net957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout958 (.A(net959),
    .X(net958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout959 (.A(net299),
    .X(net959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout961 (.A(net962),
    .X(net961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout962 (.A(net477),
    .X(net962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout963 (.A(net965),
    .X(net963),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout964 (.A(net965),
    .X(net964),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout965 (.A(net528),
    .X(net965),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout966 (.A(net967),
    .X(net966),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout967 (.A(net522),
    .X(net967),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout968 (.A(net969),
    .X(net968),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout969 (.A(net970),
    .X(net969),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout970 (.A(\DP_1.matrix[40] ),
    .X(net970),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout971 (.A(net972),
    .X(net971),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout972 (.A(net491),
    .X(net972),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout973 (.A(\DP_1.matrix[38] ),
    .X(net973),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout974 (.A(net371),
    .X(net974),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout975 (.A(net412),
    .X(net975),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout976 (.A(net412),
    .X(net976),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout977 (.A(net281),
    .X(net977),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout978 (.A(net979),
    .X(net978),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout979 (.A(net980),
    .X(net979),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout980 (.A(net505),
    .X(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout981 (.A(net982),
    .X(net981),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout982 (.A(net502),
    .X(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout983 (.A(net984),
    .X(net983),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout984 (.A(net503),
    .X(net984),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout985 (.A(net986),
    .X(net985),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout986 (.A(net510),
    .X(net986),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout987 (.A(net988),
    .X(net987),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout988 (.A(net509),
    .X(net988),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout989 (.A(net402),
    .X(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout990 (.A(\DP_1.matrix[2] ),
    .X(net990),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout991 (.A(net392),
    .X(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout992 (.A(\DP_1.matrix[1] ),
    .X(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout993 (.A(net358),
    .X(net993),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout994 (.A(\DP_4.matrix[80] ),
    .X(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout995 (.A(\DP_4.matrix[44] ),
    .X(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout996 (.A(net476),
    .X(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout997 (.A(net316),
    .X(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout998 (.A(\DP_3.matrix[80] ),
    .X(net998),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout999 (.A(net352),
    .X(net999),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1000 (.A(\DP_3.matrix[44] ),
    .X(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1001 (.A(net441),
    .X(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1002 (.A(\DP_3.matrix[8] ),
    .X(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1003 (.A(\DP_2.matrix[80] ),
    .X(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1004 (.A(net390),
    .X(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1005 (.A(net490),
    .X(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1006 (.A(net1007),
    .X(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1007 (.A(\DP_1.matrix[80] ),
    .X(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1008 (.A(net1009),
    .X(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1009 (.A(net403),
    .X(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1010 (.A(net445),
    .X(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1011 (.A(\DP_1.matrix[8] ),
    .X(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1012 (.A(net1013),
    .X(net1012),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1013 (.A(net1016),
    .X(net1013),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1014 (.A(net1016),
    .X(net1014),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1015 (.A(net1016),
    .X(net1015),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1016 (.A(net1025),
    .X(net1016),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1017 (.A(net1021),
    .X(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1018 (.A(net1021),
    .X(net1018),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1019 (.A(net1020),
    .X(net1019),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1020 (.A(net1021),
    .X(net1020),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1021 (.A(net1025),
    .X(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1022 (.A(net1023),
    .X(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1023 (.A(net1024),
    .X(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1024 (.A(net1025),
    .X(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1025 (.A(net1098),
    .X(net1025),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1026 (.A(net1030),
    .X(net1026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1027 (.A(net1030),
    .X(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1028 (.A(net1030),
    .X(net1028),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1029 (.A(net1030),
    .X(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1030 (.A(net1038),
    .X(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1031 (.A(net1034),
    .X(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1032 (.A(net1034),
    .X(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1033 (.A(net1034),
    .X(net1033),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1034 (.A(net1038),
    .X(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1035 (.A(net1037),
    .X(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1036 (.A(net1037),
    .X(net1036),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1037 (.A(net1038),
    .X(net1037),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1038 (.A(net1098),
    .X(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1039 (.A(net1040),
    .X(net1039),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1040 (.A(net1042),
    .X(net1040),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1041 (.A(net1042),
    .X(net1041),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1042 (.A(net1063),
    .X(net1042),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1043 (.A(net1044),
    .X(net1043),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1044 (.A(net1045),
    .X(net1044),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1045 (.A(net1048),
    .X(net1045),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1046 (.A(net1047),
    .X(net1046),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1047 (.A(net1048),
    .X(net1047),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1048 (.A(net1063),
    .X(net1048),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1049 (.A(net1053),
    .X(net1049),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1050 (.A(net1053),
    .X(net1050),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1051 (.A(net1053),
    .X(net1051),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1052 (.A(net1053),
    .X(net1052),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1053 (.A(net1063),
    .X(net1053),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1054 (.A(net1056),
    .X(net1054),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1055 (.A(net1056),
    .X(net1055),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1056 (.A(net1063),
    .X(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1057 (.A(net1058),
    .X(net1057),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1058 (.A(net1059),
    .X(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1059 (.A(net1062),
    .X(net1059),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1060 (.A(net1062),
    .X(net1060),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1061 (.A(net1062),
    .X(net1061),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1062 (.A(net1063),
    .X(net1062),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1063 (.A(net1098),
    .X(net1063),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1064 (.A(net1066),
    .X(net1064),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1065 (.A(net1066),
    .X(net1065),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1066 (.A(net1077),
    .X(net1066),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1067 (.A(net1069),
    .X(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1068 (.A(net1069),
    .X(net1068),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1069 (.A(net1071),
    .X(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1070 (.A(net1071),
    .X(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1071 (.A(net1077),
    .X(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1072 (.A(net1074),
    .X(net1072),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1073 (.A(net1074),
    .X(net1073),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1074 (.A(net1075),
    .X(net1074),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1075 (.A(net1077),
    .X(net1075),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1076 (.A(net1077),
    .X(net1076),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1077 (.A(net1098),
    .X(net1077),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1078 (.A(net1079),
    .X(net1078),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1079 (.A(net1087),
    .X(net1079),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1080 (.A(net1082),
    .X(net1080),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1081 (.A(net1082),
    .X(net1081),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1082 (.A(net1087),
    .X(net1082),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1083 (.A(net1084),
    .X(net1083),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1084 (.A(net1087),
    .X(net1084),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1085 (.A(net1086),
    .X(net1085),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1086 (.A(net1087),
    .X(net1086),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1087 (.A(net1098),
    .X(net1087),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1088 (.A(net1091),
    .X(net1088),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1089 (.A(net1090),
    .X(net1089),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1090 (.A(net1091),
    .X(net1090),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1091 (.A(net1097),
    .X(net1091),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1092 (.A(net1095),
    .X(net1092),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1093 (.A(net1094),
    .X(net1093),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1094 (.A(net1095),
    .X(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1095 (.A(net1097),
    .X(net1095),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1096 (.A(net1097),
    .X(net1096),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1097 (.A(net1098),
    .X(net1097),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1098 (.A(rst_n),
    .X(net1098),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi heichips25_SDR_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_41_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_45_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_46_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_50_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_51_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_52_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_54_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_55_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_56_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_57_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_58_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_59_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_60_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_61_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_62_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_63_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_64_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_65_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_66_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload0 (.A(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload3 (.A(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload4 (.A(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload5 (.A(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload6 (.A(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload7 (.A(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload8 (.A(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload9 (.A(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload10 (.A(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload11 (.A(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload12 (.A(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload13 (.VDD(VPWR),
    .A(clknet_leaf_65_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload14 (.VDD(VPWR),
    .A(clknet_leaf_66_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload15 (.VDD(VPWR),
    .A(clknet_leaf_28_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload16 (.VDD(VPWR),
    .A(clknet_leaf_27_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_56_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_57_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_59_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload21 (.VDD(VPWR),
    .A(clknet_leaf_50_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload23 (.VDD(VPWR),
    .A(clknet_leaf_33_clk),
    .VSS(VGND));
 sg13g2_inv_8 clkload24 (.A(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac1.sum_lvl1_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac2.sum_lvl1_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac1.products_ff[144] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac1.products_ff[149] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac2.products_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac1.sum_lvl1_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac2.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac2.sum_lvl2_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac1.sum_lvl1_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac2.sum_lvl1_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac1.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac2.sum_lvl1_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac1.sum_lvl2_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mac2.products_ff[145] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mac1.sum_lvl2_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mac2.sum_lvl2_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mac1.products_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mac1.sum_lvl2_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mac2.sum_lvl1_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mac1.products_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mac1.products_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mac2.products_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mac2.sum_lvl1_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mac1.products_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mac1.products_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mac2.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mac2.sum_lvl2_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mac1.products_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mac2.sum_lvl1_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mac1.sum_lvl2_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mac1.sum_lvl1_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mac2.sum_lvl1_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mac2.sum_lvl1_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mac1.sum_lvl2_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mac1.products_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mac1.products_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mac2.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mac2.products_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mac2.products_ff[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mac1.products_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mac1.sum_lvl1_ff[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mac2.sum_lvl2_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mac2.sum_lvl2_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mac2.sum_lvl1_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mac2.sum_lvl2_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mac1.products_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mac1.sum_lvl1_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mac2.sum_lvl1_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mac1.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mac2.sum_lvl1_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mac2.sum_lvl1_ff[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mac1.products_ff[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mac2.products_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mac1.sum_lvl1_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mac2.sum_lvl1_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mac1.sum_lvl1_ff[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac2.products_ff[148] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mac1.products_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac1.products_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mac1.sum_lvl1_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac1.sum_lvl1_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mac1.products_ff[151] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac1.sum_lvl1_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mac2.sum_lvl1_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac2.sum_lvl1_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mac1.sum_lvl2_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mac2.sum_lvl1_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mac2.sum_lvl1_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mac2.sum_lvl1_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mac1.sum_lvl1_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mac2.products_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mac2.products_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mac2.sum_lvl2_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mac1.sum_lvl1_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mac1.sum_lvl1_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mac1.sum_lvl1_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mac2.sum_lvl2_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mac2.sum_lvl1_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mac2.sum_lvl1_ff[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mac1.sum_lvl2_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mac2.products_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mac2.products_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mac1.sum_lvl2_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mac2.sum_lvl1_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mac2.sum_lvl1_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mac1.sum_lvl1_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mac1.sum_lvl1_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mac2.sum_lvl1_ff[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mac1.sum_lvl2_ff[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mac2.sum_lvl1_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mac1.sum_lvl1_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mac2.products_ff[144] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mac2.sum_lvl1_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mac1.products_ff[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac1.sum_lvl1_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mac1.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac2.sum_lvl2_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mac2.products_ff[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mac2.sum_lvl1_ff[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mac2.sum_lvl1_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mac2.sum_lvl1_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac1.sum_lvl2_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mac1.sum_lvl2_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mac1.products_ff[142] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mac2.sum_lvl2_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mac1.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mac1.products_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mac1.sum_lvl1_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mac1.products_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mac1.products_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mac1.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mac1.products_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mac1.sum_lvl1_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mac2.sum_lvl1_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mac2.sum_lvl1_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mac2.sum_lvl1_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac1.sum_lvl1_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mac1.sum_lvl2_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mac2.sum_lvl1_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac1.sum_lvl1_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mac1.products_ff[139] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mac1.sum_lvl1_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac2.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mac1.sum_lvl1_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mac2.products_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mac1.products_ff[143] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mac2.products_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mac2.products_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mac2.sum_lvl2_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mac1.sum_lvl1_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mac1.sum_lvl2_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac1.sum_lvl1_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mac1.sum_lvl1_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mac2.sum_lvl2_ff[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mac1.products_ff[141] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mac1.products_ff[147] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mac1.products_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mac2.sum_lvl1_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mac1.products_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mac1.sum_lvl1_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac1.sum_lvl2_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mac2.sum_lvl1_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mac1.sum_lvl1_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mac2.products_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mac2.products_ff[141] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mac2.products_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mac1.sum_lvl1_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mac2.sum_lvl1_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mac2.products_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mac2.sum_lvl1_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac2.products_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mac1.sum_lvl1_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mac1.sum_lvl1_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mac2.sum_lvl1_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mac2.products_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mac2.sum_lvl1_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mac1.sum_lvl1_ff[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mac1.products_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mac2.products_ff[151] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mac2.sum_lvl1_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mac1.sum_lvl1_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mac1.products_ff[148] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mac2.products_ff[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mac1.products_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mac1.sum_lvl1_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mac1.products_ff[150] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mac1.sum_lvl1_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mac2.products_ff[143] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mac2.products_ff[147] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mac1.products_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mac2.products_ff[146] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mac1.products_ff[140] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mac1.sum_lvl1_ff[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mac2.products_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mac1.sum_lvl1_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mac1.sum_lvl1_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mac1.sum_lvl1_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mac2.products_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mac2.products_ff[149] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mac1.sum_lvl1_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mac1.sum_lvl1_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mac2.sum_lvl1_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mac2.products_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mac1.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mac1.products_ff[146] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mac1.sum_lvl2_ff[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mac2.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mac2.products_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mac2.products_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mac1.products_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mac1.products_ff[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mac1.products_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mac2.sum_lvl2_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mac2.products_ff[139] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mac2.sum_lvl1_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mac1.sum_lvl1_ff[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mac1.products_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold198 (.A(\mac2.sum_lvl1_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mac1.sum_lvl1_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mac1.products_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mac2.sum_lvl2_ff[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold202 (.A(\mac1.sum_lvl1_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mac2.sum_lvl1_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mac2.sum_lvl1_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold205 (.A(\mac2.products_ff[142] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mac2.sum_lvl1_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mac1.products_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mac2.products_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mac1.products_ff[138] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mac2.sum_lvl1_ff[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mac2.sum_lvl2_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mac2.products_ff[138] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mac2.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mac2.products_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mac2.products_ff[140] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mac2.sum_lvl2_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mac1.products_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mac2.products_ff[150] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mac1.products_ff[145] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mac1.sum_lvl2_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mac2.products_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mac2.products_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mac2.products_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mac2.products_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mac1.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mac2.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold229 (.A(\DP_1.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold230 (.A(\DP_1.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold231 (.A(\DP_3.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold232 (.A(\DP_4.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold233 (.A(\DP_4.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold234 (.A(\DP_3.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold235 (.A(\DP_2.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold236 (.A(\DP_1.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold237 (.A(\DP_2.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold238 (.A(\DP_1.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold239 (.A(\DP_3.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold240 (.A(\DP_2.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold241 (.A(\DP_1.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold242 (.A(\DP_4.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold243 (.A(\mac1.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold245 (.A(\mac1.sum_lvl2_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold246 (.A(_2138_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold248 (.A(\DP_4.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1717_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold251 (.A(\mac2.sum_lvl2_ff[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0039_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold253 (.A(\mac1.sum_lvl3_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold254 (.A(_2170_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold256 (.A(\DP_4.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold257 (.A(\DP_1.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold258 (.A(\DP_3.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold259 (.A(\DP_1.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold260 (.A(\DP_4.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold261 (.A(\DP_2.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold262 (.A(\DP_3.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold263 (.A(\DP_4.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold264 (.A(\DP_1.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mac2.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0048_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold267 (.A(\DP_2.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold268 (.A(\DP_3.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold269 (.A(\DP_4.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold270 (.A(\DP_2.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold271 (.A(\mac2.sum_lvl3_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold272 (.A(_2293_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0051_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold274 (.A(\DP_4.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold275 (.A(\DP_4.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold276 (.A(\DP_3.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mac1.sum_lvl3_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold278 (.A(_2154_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mac2.sum_lvl2_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold281 (.A(_2200_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0040_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mac1.sum_lvl3_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold284 (.A(_2183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold286 (.A(\DP_1.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold287 (.A(\DP_3.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold288 (.A(\DP_4.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold289 (.A(\DP_3.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold290 (.A(\DP_4.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold291 (.A(\DP_4.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold292 (.A(\mac1.sum_lvl2_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold293 (.A(_2087_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold295 (.A(\DP_2.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold296 (.A(\DP_1.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold297 (.A(\DP_4.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold298 (.A(\mac2.sum_lvl3_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold299 (.A(_2279_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0063_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold301 (.A(\mac1.sum_lvl3_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold302 (.A(_2187_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold304 (.A(\DP_4.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold305 (.A(\DP_2.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold306 (.A(\DP_2.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mac2.sum_lvl3_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold308 (.A(_2301_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold310 (.A(\DP_4.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0247_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold312 (.A(\DP_3.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold313 (.A(\mac1.sum_lvl3_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold314 (.A(_2151_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold316 (.A(\DP_4.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold317 (.A(\DP_2.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold318 (.A(\DP_1.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold319 (.A(\DP_4.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold320 (.A(\mac2.sum_lvl2_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold321 (.A(_2203_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0041_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold323 (.A(\DP_3.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold324 (.A(\DP_3.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold325 (.A(\DP_3.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold326 (.A(\DP_4.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold327 (.A(\mac2.sum_lvl3_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold328 (.A(_2303_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold330 (.A(\DP_3.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold331 (.A(\DP_1.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold332 (.A(\DP_3.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold333 (.A(\mac1.sum_lvl3_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold334 (.A(_2190_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold336 (.A(\DP_4.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold337 (.A(\mac1.sum_lvl3_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold338 (.A(_2173_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold340 (.A(\mac2.sum_lvl3_ff[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold341 (.A(_2281_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold343 (.A(\mac1.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold344 (.A(_2148_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold346 (.A(\DP_3.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold347 (.A(\DP_2.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold348 (.A(\DP_2.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0198_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold350 (.A(\DP_2.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold351 (.A(\DP_2.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold352 (.A(\DP_1.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold353 (.A(\mac1.sum_lvl3_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold354 (.A(_2176_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold356 (.A(\DP_3.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold357 (.A(_2571_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold358 (.A(\mac2.sum_lvl3_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold359 (.A(_2295_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold360 (.A(_2296_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0052_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold362 (.A(\DP_1.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold363 (.A(\DP_1.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold364 (.A(\DP_4.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold365 (.A(\mac1.sum_lvl3_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold366 (.A(_2164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold367 (.A(_2165_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold369 (.A(\mac1.sum_lvl3_ff[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold370 (.A(_2193_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold372 (.A(\DP_1.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold373 (.A(\DP_4.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold374 (.A(\DP_2.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold375 (.A(\mac1.sum_lvl2_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold376 (.A(_2090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold378 (.A(\mac2.sum_lvl3_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold379 (.A(_2264_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0059_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold381 (.A(\DP_3.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold382 (.A(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold383 (.A(\mac2.sum_lvl3_ff[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold384 (.A(_2284_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold385 (.A(_2286_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold387 (.A(\DP_2.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold388 (.A(\DP_4.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold389 (.A(\mac1.sum_lvl3_ff[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold391 (.A(\DP_2.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold392 (.A(_2551_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold393 (.A(\mac1.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold394 (.A(_2145_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold396 (.A(\mac2.sum_lvl3_ff[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold397 (.A(_2270_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold398 (.A(_2276_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold400 (.A(\DP_4.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold401 (.A(\DP_3.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold402 (.A(\DP_2.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold403 (.A(\DP_2.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold404 (.A(\DP_2.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold405 (.A(\DP_1.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0160_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold407 (.A(\DP_3.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold408 (.A(\mac2.sum_lvl2_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold409 (.A(_2209_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold411 (.A(\mac2.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold412 (.A(_2255_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold414 (.A(\mac2.sum_lvl3_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold415 (.A(_2261_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0058_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold417 (.A(\mac2.sum_lvl3_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold418 (.A(_2266_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold419 (.A(_2269_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0060_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold421 (.A(\mac2.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold422 (.A(_2206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold424 (.A(\DP_2.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold425 (.A(\DP_4.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold426 (.A(\DP_2.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold427 (.A(\DP_4.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold428 (.A(\mac1.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold429 (.A(_2136_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold431 (.A(\DP_2.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold432 (.A(\DP_3.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold433 (.A(\DP_3.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold434 (.A(\mac2.sum_lvl3_ff[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold436 (.A(\DP_4.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold437 (.A(\DP_1.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold438 (.A(\mac1.sum_lvl2_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold439 (.A(_2130_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold440 (.A(_2131_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold442 (.A(\DP_4.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold443 (.A(\mac1.sum_lvl3_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold444 (.A(_2156_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold445 (.A(_2159_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold447 (.A(\mac2.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold448 (.A(_2258_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold450 (.A(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold451 (.A(\DP_1.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold452 (.A(\DP_3.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold453 (.A(\DP_3.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold454 (.A(\mac1.sum_lvl2_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold455 (.A(_2093_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold457 (.A(\DP_3.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold458 (.A(\DP_3.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold459 (.A(\mac1.sum_lvl2_ff[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold460 (.A(_2105_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold462 (.A(\DP_1.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold463 (.A(\DP_1.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold464 (.A(\DP_2.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold465 (.A(\DP_1.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold466 (.A(\mac2.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold467 (.A(_2215_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold469 (.A(\DP_1.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold470 (.A(\DP_1.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold471 (.A(\mac2.sum_lvl2_ff[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold472 (.A(_2237_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0036_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold474 (.A(\mac1.sum_lvl2_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold475 (.A(_2101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold476 (.A(_2104_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold477 (.A(\DP_3.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold478 (.A(\mac1.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold479 (.A(_2161_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold480 (.A(_2162_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold482 (.A(\DP_1.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold483 (.A(\DP_2.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold484 (.A(\mac2.sum_lvl2_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold485 (.A(_2211_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold486 (.A(_2214_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold488 (.A(\DP_1.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold489 (.A(\mac1.sum_lvl2_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold490 (.A(_2099_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold491 (.A(\mac2.sum_lvl2_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold492 (.A(_2248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold493 (.A(\mac1.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold494 (.A(_2096_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold495 (.A(\mac1.sum_lvl2_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold496 (.A(_2128_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold497 (.A(\mac1.sum_lvl2_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold498 (.A(_2116_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold499 (.A(\mac2.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold500 (.A(_2273_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold502 (.A(\mac2.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold503 (.A(_2224_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold504 (.A(\mac2.sum_lvl2_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold505 (.A(_2226_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold506 (.A(\mac1.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold507 (.A(_2114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold508 (.A(\mac1.sum_lvl2_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net548));
 sg13g2_fill_2 FILLER_0_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net33;
 assign uio_oe[1] = net34;
 assign uio_oe[2] = net35;
 assign uio_oe[3] = net36;
 assign uio_oe[4] = net37;
 assign uio_oe[5] = net38;
 assign uio_oe[6] = net39;
 assign uio_oe[7] = net40;
endmodule
