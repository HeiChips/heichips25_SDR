* NGSPICE file created from heichips25_SDR.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

.subckt heichips25_SDR VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ _2747_ net947 net894 net892 net950 VPWR VGND sg13g2_a22oi_1
X_3086_ _2675_ VPWR _2680_ VGND _2676_ _2678_ sg13g2_o21ai_1
XFILLER_36_962 VPWR VGND sg13g2_decap_8
XFILLER_23_601 VPWR VGND sg13g2_decap_8
X_3988_ VGND VPWR _0788_ _0791_ _0832_ _0831_ sg13g2_a21oi_1
X_5727_ _2430_ _2434_ _2435_ VPWR VGND sg13g2_nor2b_1
X_5658_ DP_1.Q_range.out_data\[3\] DP_1.I_range.out_data\[3\] _2367_ VPWR VGND sg13g2_xor2_1
X_5589_ _2312_ mac1.total_sum\[3\] mac2.total_sum\[3\] VPWR VGND sg13g2_nand2_1
X_4609_ _1424_ net881 net825 VPWR VGND sg13g2_nand2_1
Xhold362 DP_1.matrix\[2\] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold351 DP_2.matrix\[36\] VPWR VGND net391 sg13g2_dlygate4sd3_1
Xhold340 mac2.sum_lvl3_ff\[30\] VPWR VGND net380 sg13g2_dlygate4sd3_1
Xhold373 DP_4.matrix\[6\] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold395 _0024_ VPWR VGND net435 sg13g2_dlygate4sd3_1
XFILLER_2_549 VPWR VGND sg13g2_fill_2
Xhold384 _2284_ VPWR VGND net424 sg13g2_dlygate4sd3_1
Xfanout820 net428 net820 VPWR VGND sg13g2_buf_8
Xfanout842 net843 net842 VPWR VGND sg13g2_buf_1
Xfanout831 net832 net831 VPWR VGND sg13g2_buf_2
Xfanout875 DP_3.matrix\[6\] net875 VPWR VGND sg13g2_buf_8
Xfanout853 net372 net853 VPWR VGND sg13g2_buf_1
Xfanout864 net492 net864 VPWR VGND sg13g2_buf_8
Xfanout897 net310 net897 VPWR VGND sg13g2_buf_2
Xfanout886 net365 net886 VPWR VGND sg13g2_buf_8
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_33_409 VPWR VGND sg13g2_fill_2
XFILLER_42_910 VPWR VGND sg13g2_decap_8
XFILLER_42_987 VPWR VGND sg13g2_decap_8
XFILLER_6_877 VPWR VGND sg13g2_fill_1
XFILLER_3_56 VPWR VGND sg13g2_fill_1
XFILLER_49_553 VPWR VGND sg13g2_fill_1
XFILLER_49_586 VPWR VGND sg13g2_decap_8
XFILLER_18_962 VPWR VGND sg13g2_decap_8
XFILLER_17_461 VPWR VGND sg13g2_fill_1
X_4960_ _1760_ net850 net789 VPWR VGND sg13g2_nand2_1
X_4891_ _1698_ _1697_ _1694_ VPWR VGND sg13g2_nand2b_1
X_3911_ _0756_ net974 net908 VPWR VGND sg13g2_nand2_1
XFILLER_32_420 VPWR VGND sg13g2_fill_1
XFILLER_33_965 VPWR VGND sg13g2_decap_8
X_3842_ _0689_ net972 net912 VPWR VGND sg13g2_nand2_1
XFILLER_20_637 VPWR VGND sg13g2_decap_4
XFILLER_32_497 VPWR VGND sg13g2_fill_1
XFILLER_9_671 VPWR VGND sg13g2_fill_2
X_3773_ VGND VPWR _0616_ _0619_ _0623_ _0617_ sg13g2_a21oi_1
X_5512_ _0055_ _2249_ _2252_ VPWR VGND sg13g2_xnor2_1
X_6492_ net1026 VGND VPWR net8 DP_1.Q_range.out_data\[6\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5443_ mac2.sum_lvl2_ff\[21\] net320 _2199_ VPWR VGND sg13g2_and2_1
X_5374_ net434 _2143_ _0024_ VPWR VGND sg13g2_xor2_1
X_4325_ _1129_ VPWR _1154_ VGND _1150_ _1152_ sg13g2_o21ai_1
X_4256_ _1083_ _1085_ _1086_ VPWR VGND sg13g2_nor2b_1
X_3207_ _2798_ net896 net1006 VPWR VGND sg13g2_nand2_1
X_4187_ _1018_ _1017_ _1020_ VPWR VGND sg13g2_xor2_1
X_3138_ _2731_ _2729_ _2730_ VPWR VGND sg13g2_nand2_1
X_3069_ _2640_ VPWR _2663_ VGND _2617_ _2638_ sg13g2_o21ai_1
Xhold170 mac1.products_ff\[81\] VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold181 mac1.sum_lvl1_ff\[47\] VPWR VGND net221 sg13g2_dlygate4sd3_1
Xhold192 mac1.products_ff\[80\] VPWR VGND net232 sg13g2_dlygate4sd3_1
XFILLER_37_95 VPWR VGND sg13g2_fill_2
XFILLER_42_740 VPWR VGND sg13g2_fill_2
XFILLER_14_431 VPWR VGND sg13g2_fill_2
XFILLER_18_1004 VPWR VGND sg13g2_decap_8
XFILLER_14_442 VPWR VGND sg13g2_fill_2
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_30_913 VPWR VGND sg13g2_decap_8
XFILLER_6_652 VPWR VGND sg13g2_fill_1
XFILLER_6_674 VPWR VGND sg13g2_fill_1
X_4110_ _0950_ _0932_ _0949_ VPWR VGND sg13g2_nand2_1
XFILLER_25_1008 VPWR VGND sg13g2_decap_8
X_5090_ _1884_ _1885_ _1866_ _1887_ VPWR VGND sg13g2_nand3_1
X_4041_ VGND VPWR _0883_ _0856_ _0854_ sg13g2_or2_1
X_5992_ net1043 VGND VPWR _0070_ mac1.products_ff\[1\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_4943_ net799 net795 net849 net847 _1744_ VPWR VGND sg13g2_and4_1
X_4874_ _1682_ _1652_ _1680_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_401 VPWR VGND sg13g2_fill_1
X_3825_ _0661_ VPWR _0673_ VGND _0669_ _0671_ sg13g2_o21ai_1
X_3756_ _0609_ _0592_ _0610_ VPWR VGND sg13g2_xor2_1
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
X_6475_ net1012 VGND VPWR net489 mac2.total_sum\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_5426_ _2187_ mac1.sum_lvl3_ff\[33\] net341 VPWR VGND sg13g2_xnor2_1
X_3687_ _0544_ net982 DP_2.matrix\[7\] VPWR VGND sg13g2_nand2_1
X_5357_ VGND VPWR mac1.sum_lvl2_ff\[32\] mac1.sum_lvl2_ff\[13\] _2133_ _2131_ sg13g2_a21oi_1
X_5288_ _2065_ VPWR _2078_ VGND _2039_ _2063_ sg13g2_o21ai_1
X_4308_ _1137_ _1136_ _1135_ VPWR VGND sg13g2_nand2b_1
X_4239_ _1067_ _1066_ _1061_ _1070_ VPWR VGND sg13g2_a21o_1
XFILLER_16_729 VPWR VGND sg13g2_fill_1
XFILLER_8_906 VPWR VGND sg13g2_fill_1
XFILLER_12_957 VPWR VGND sg13g2_decap_8
XFILLER_23_53 VPWR VGND sg13g2_fill_1
XFILLER_3_600 VPWR VGND sg13g2_fill_2
XFILLER_38_309 VPWR VGND sg13g2_fill_2
XFILLER_47_876 VPWR VGND sg13g2_decap_8
X_3610_ _0470_ _0426_ _0429_ VPWR VGND sg13g2_nand2_1
X_4590_ _1395_ _1403_ _1405_ _1406_ VPWR VGND sg13g2_or3_1
XFILLER_7_950 VPWR VGND sg13g2_decap_8
X_3541_ _0402_ _0356_ _0399_ VPWR VGND sg13g2_xnor2_1
X_3472_ _0332_ _0331_ _0326_ _0335_ VPWR VGND sg13g2_a21o_1
X_6260_ net1052 VGND VPWR net66 mac2.sum_lvl1_ff\[73\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6191_ net1085 VGND VPWR net94 mac1.sum_lvl2_ff\[12\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5211_ VGND VPWR _1972_ _1975_ _2005_ _1970_ sg13g2_a21oi_1
X_5142_ _1938_ _1891_ _1894_ _1935_ VPWR VGND sg13g2_and3_1
X_5073_ VGND VPWR _1870_ _1868_ _1827_ sg13g2_or2_1
XFILLER_49_180 VPWR VGND sg13g2_fill_2
X_4024_ VGND VPWR _0828_ _0830_ _0867_ _0866_ sg13g2_a21oi_1
XFILLER_37_331 VPWR VGND sg13g2_fill_2
XFILLER_38_865 VPWR VGND sg13g2_decap_8
XFILLER_25_526 VPWR VGND sg13g2_fill_2
X_5975_ net805 _0257_ VPWR VGND sg13g2_buf_1
XFILLER_21_721 VPWR VGND sg13g2_fill_1
X_4926_ DP_4.matrix\[73\] net851 net799 _1728_ VPWR VGND net848 sg13g2_nand4_1
X_4857_ _1666_ _1661_ _1665_ VPWR VGND sg13g2_nand2_1
X_3808_ _0656_ net977 net911 VPWR VGND sg13g2_nand2_1
X_4788_ _1599_ _1571_ _1598_ VPWR VGND sg13g2_nand2_1
X_3739_ _0593_ _0569_ _0594_ VPWR VGND sg13g2_xor2_1
X_6458_ net1058 VGND VPWR net322 mac2.sum_lvl3_ff\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5409_ _2173_ mac1.sum_lvl3_ff\[30\] net377 VPWR VGND sg13g2_xnor2_1
X_6389_ net1059 VGND VPWR net223 mac2.sum_lvl1_ff\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_44_879 VPWR VGND sg13g2_decap_8
XFILLER_31_507 VPWR VGND sg13g2_fill_2
XFILLER_43_389 VPWR VGND sg13g2_fill_1
XFILLER_43_378 VPWR VGND sg13g2_fill_1
XFILLER_4_975 VPWR VGND sg13g2_decap_8
XFILLER_3_485 VPWR VGND sg13g2_fill_1
XFILLER_3_474 VPWR VGND sg13g2_fill_2
XFILLER_35_802 VPWR VGND sg13g2_fill_2
XFILLER_46_172 VPWR VGND sg13g2_fill_1
XFILLER_34_312 VPWR VGND sg13g2_fill_1
XFILLER_15_570 VPWR VGND sg13g2_fill_2
X_5760_ _2464_ _2465_ _2466_ _2467_ VPWR VGND sg13g2_nor3_1
X_5691_ _2395_ _2399_ _2400_ VPWR VGND sg13g2_nor2b_1
XFILLER_15_592 VPWR VGND sg13g2_fill_2
X_4711_ _1523_ _1522_ _1454_ _1524_ VPWR VGND sg13g2_a21o_1
XFILLER_30_573 VPWR VGND sg13g2_fill_2
X_4642_ _1437_ _1427_ _1435_ _1456_ VPWR VGND sg13g2_a21o_1
X_4573_ _1381_ VPWR _1389_ VGND _1373_ _1383_ sg13g2_o21ai_1
X_3524_ _0374_ VPWR _0385_ VGND _0353_ _0375_ sg13g2_o21ai_1
X_6312_ net1049 VGND VPWR net251 mac2.sum_lvl3_ff\[25\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3455_ _0316_ _0315_ _0318_ VPWR VGND sg13g2_xor2_1
X_6243_ net1039 VGND VPWR net136 mac1.sum_lvl1_ff\[72\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3386_ _2968_ _2961_ _2967_ VPWR VGND sg13g2_nand2_1
X_6174_ net1084 VGND VPWR net257 mac1.sum_lvl1_ff\[47\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5125_ _1877_ VPWR _1921_ VGND _1875_ _1878_ sg13g2_o21ai_1
X_5056_ _1854_ _1852_ _1853_ VPWR VGND sg13g2_nand2_1
XFILLER_38_640 VPWR VGND sg13g2_fill_1
X_4007_ _0822_ VPWR _0850_ VGND _0816_ _0823_ sg13g2_o21ai_1
XFILLER_38_695 VPWR VGND sg13g2_decap_4
X_5958_ net863 _0232_ VPWR VGND sg13g2_buf_1
X_4909_ _1715_ _1709_ _1714_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_359 VPWR VGND sg13g2_fill_2
X_5889_ _2571_ net873 net762 VPWR VGND sg13g2_nand2_1
XFILLER_1_934 VPWR VGND sg13g2_decap_8
XFILLER_49_905 VPWR VGND sg13g2_decap_8
Xhold30 mac1.sum_lvl2_ff\[39\] VPWR VGND net70 sg13g2_dlygate4sd3_1
Xhold41 mac1.sum_lvl1_ff\[86\] VPWR VGND net81 sg13g2_dlygate4sd3_1
Xhold74 mac1.sum_lvl1_ff\[2\] VPWR VGND net114 sg13g2_dlygate4sd3_1
Xhold52 mac1.products_ff\[69\] VPWR VGND net92 sg13g2_dlygate4sd3_1
XFILLER_21_1011 VPWR VGND sg13g2_decap_8
Xhold63 mac1.sum_lvl1_ff\[14\] VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold96 mac1.products_ff\[136\] VPWR VGND net136 sg13g2_dlygate4sd3_1
XFILLER_28_150 VPWR VGND sg13g2_fill_2
Xhold85 mac2.sum_lvl1_ff\[45\] VPWR VGND net125 sg13g2_dlygate4sd3_1
XFILLER_44_643 VPWR VGND sg13g2_fill_1
XFILLER_16_334 VPWR VGND sg13g2_fill_2
XFILLER_45_84 VPWR VGND sg13g2_fill_2
XFILLER_43_175 VPWR VGND sg13g2_fill_2
XFILLER_12_551 VPWR VGND sg13g2_fill_2
XFILLER_40_871 VPWR VGND sg13g2_decap_8
XFILLER_8_599 VPWR VGND sg13g2_decap_4
XFILLER_4_761 VPWR VGND sg13g2_fill_2
X_3240_ _2802_ VPWR _2830_ VGND _2796_ _2803_ sg13g2_o21ai_1
X_3171_ _2763_ _2743_ _2761_ _2762_ VPWR VGND sg13g2_and3_1
Xfanout1050 net1053 net1050 VPWR VGND sg13g2_buf_8
Xfanout1083 net1084 net1083 VPWR VGND sg13g2_buf_8
Xfanout1072 net1074 net1072 VPWR VGND sg13g2_buf_8
XFILLER_39_459 VPWR VGND sg13g2_fill_2
Xfanout1061 net1062 net1061 VPWR VGND sg13g2_buf_8
XFILLER_48_982 VPWR VGND sg13g2_decap_8
Xfanout1094 net1095 net1094 VPWR VGND sg13g2_buf_8
X_5812_ net804 net779 _2518_ VPWR VGND sg13g2_nor2_1
X_5743_ net768 VPWR _2450_ VGND net1001 net777 sg13g2_o21ai_1
XFILLER_16_890 VPWR VGND sg13g2_fill_1
XFILLER_31_871 VPWR VGND sg13g2_decap_8
X_5674_ net977 net993 net774 _2383_ VPWR VGND sg13g2_mux2_1
X_4625_ _1438_ _1439_ _1421_ _1440_ VPWR VGND sg13g2_nand3_1
Xhold500 _2273_ VPWR VGND net540 sg13g2_dlygate4sd3_1
X_4556_ VGND VPWR _1373_ _1372_ _1370_ sg13g2_or2_1
X_3507_ _0366_ _0367_ _0361_ _0369_ VPWR VGND sg13g2_nand3_1
X_4487_ _1271_ _1310_ _1311_ VPWR VGND sg13g2_nor2_1
X_3438_ _0299_ _0300_ _0294_ _0302_ VPWR VGND sg13g2_nand3_1
X_6226_ net1065 VGND VPWR net213 mac1.sum_lvl2_ff\[53\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_6157_ net1054 VGND VPWR _0262_ DP_4.matrix\[74\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3369_ VGND VPWR _2924_ _2947_ _2954_ _2949_ sg13g2_a21oi_1
X_5108_ _1904_ net852 net994 VPWR VGND sg13g2_nand2_1
X_6088_ net1025 VGND VPWR _0098_ mac1.products_ff\[149\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_39_993 VPWR VGND sg13g2_decap_8
X_5039_ _1832_ VPWR _1837_ VGND _1833_ _1835_ sg13g2_o21ai_1
XFILLER_26_676 VPWR VGND sg13g2_decap_8
Xoutput31 net31 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_49_757 VPWR VGND sg13g2_decap_8
XFILLER_0_274 VPWR VGND sg13g2_fill_2
XFILLER_36_407 VPWR VGND sg13g2_fill_1
XFILLER_45_930 VPWR VGND sg13g2_decap_8
XFILLER_32_624 VPWR VGND sg13g2_fill_2
XFILLER_9_897 VPWR VGND sg13g2_fill_1
XFILLER_12_392 VPWR VGND sg13g2_fill_2
X_4410_ _1117_ _1162_ _1116_ _1237_ VPWR VGND _1202_ sg13g2_nand4_1
X_5390_ _2153_ net484 _2157_ _2158_ VPWR VGND sg13g2_nor3_1
X_4341_ _1169_ net866 net801 VPWR VGND sg13g2_nand2_1
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_4272_ _1102_ _1095_ _1100_ _1101_ VPWR VGND sg13g2_and3_1
X_6011_ net1067 VGND VPWR _0078_ mac1.products_ff\[72\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3223_ _2814_ _2768_ _2771_ _2811_ VPWR VGND sg13g2_and3_1
X_3154_ net894 net950 net892 net946 _2746_ VPWR VGND sg13g2_and4_1
X_3085_ _2675_ _2676_ _2678_ _2679_ VPWR VGND sg13g2_or3_1
XFILLER_36_941 VPWR VGND sg13g2_decap_8
X_3987_ _0829_ _0797_ _0831_ VPWR VGND sg13g2_xor2_1
X_5726_ _2431_ VPWR _2434_ VGND _2432_ _2433_ sg13g2_o21ai_1
X_5657_ VGND VPWR _2365_ _2366_ _2361_ _2360_ sg13g2_a21oi_2
X_5588_ VGND VPWR _2308_ _2310_ _2311_ _2309_ sg13g2_a21oi_1
X_4608_ _1423_ net881 net823 VPWR VGND sg13g2_nand2_1
Xhold352 DP_1.matrix\[1\] VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold341 _2281_ VPWR VGND net381 sg13g2_dlygate4sd3_1
X_4539_ VGND VPWR _1350_ _1353_ _1357_ _1351_ sg13g2_a21oi_1
Xhold330 DP_3.matrix\[1\] VPWR VGND net370 sg13g2_dlygate4sd3_1
Xhold374 DP_2.matrix\[6\] VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold363 DP_1.matrix\[44\] VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold396 mac2.sum_lvl3_ff\[27\] VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold385 _2286_ VPWR VGND net425 sg13g2_dlygate4sd3_1
Xfanout843 net308 net843 VPWR VGND sg13g2_buf_2
Xfanout821 net413 net821 VPWR VGND sg13g2_buf_8
X_6209_ net1084 VGND VPWR net217 mac1.sum_lvl2_ff\[33\] clknet_leaf_47_clk sg13g2_dfrbpq_2
Xfanout832 DP_4.matrix\[1\] net832 VPWR VGND sg13g2_buf_2
Xfanout810 DP_4.matrix\[39\] net810 VPWR VGND sg13g2_buf_1
Xfanout876 net364 net876 VPWR VGND sg13g2_buf_8
Xfanout854 DP_3.matrix\[72\] net854 VPWR VGND sg13g2_buf_8
Xfanout865 net866 net865 VPWR VGND sg13g2_buf_8
XFILLER_46_705 VPWR VGND sg13g2_fill_2
Xfanout898 net902 net898 VPWR VGND sg13g2_buf_2
Xfanout887 net888 net887 VPWR VGND sg13g2_buf_8
XFILLER_46_749 VPWR VGND sg13g2_fill_2
XFILLER_27_952 VPWR VGND sg13g2_decap_8
XFILLER_42_966 VPWR VGND sg13g2_decap_8
XFILLER_41_421 VPWR VGND sg13g2_fill_1
XFILLER_6_812 VPWR VGND sg13g2_fill_2
XFILLER_22_690 VPWR VGND sg13g2_fill_1
XFILLER_6_845 VPWR VGND sg13g2_fill_2
XFILLER_10_896 VPWR VGND sg13g2_fill_2
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_49_565 VPWR VGND sg13g2_fill_2
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
XFILLER_36_226 VPWR VGND sg13g2_fill_1
XFILLER_45_760 VPWR VGND sg13g2_fill_1
X_4890_ _1696_ _1671_ _1697_ VPWR VGND sg13g2_xor2_1
X_3910_ _0755_ net974 net906 VPWR VGND sg13g2_nand2_1
XFILLER_33_944 VPWR VGND sg13g2_decap_8
X_3841_ _0688_ net976 net910 VPWR VGND sg13g2_nand2_1
X_3772_ _0622_ net281 net504 VPWR VGND sg13g2_nand2_2
XFILLER_32_476 VPWR VGND sg13g2_fill_1
XFILLER_34_1010 VPWR VGND sg13g2_decap_8
X_5511_ mac2.sum_lvl3_ff\[1\] mac2.sum_lvl3_ff\[21\] _2252_ VPWR VGND sg13g2_xor2_1
XFILLER_9_683 VPWR VGND sg13g2_decap_4
X_6491_ net1026 VGND VPWR DP_1.Q_range.data_plus_4\[6\] DP_1.Q_range.out_data\[5\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5442_ _2195_ VPWR _2198_ VGND _2194_ _2196_ sg13g2_o21ai_1
X_5373_ net433 mac1.sum_lvl3_ff\[22\] _2145_ VPWR VGND sg13g2_xor2_1
X_4324_ _1129_ _1150_ _1152_ _1153_ VPWR VGND sg13g2_or3_1
X_4255_ VGND VPWR _1085_ _1084_ _1051_ sg13g2_or2_1
X_3206_ _2754_ VPWR _2797_ VGND _2752_ _2755_ sg13g2_o21ai_1
X_4186_ _1019_ _1017_ _1018_ VPWR VGND sg13g2_nand2_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
X_3137_ _2691_ VPWR _2730_ VGND _2692_ _2693_ sg13g2_o21ai_1
X_3068_ _2662_ _2654_ _2658_ VPWR VGND sg13g2_nand2_1
XFILLER_36_760 VPWR VGND sg13g2_fill_2
XFILLER_24_988 VPWR VGND sg13g2_decap_8
XFILLER_23_498 VPWR VGND sg13g2_fill_2
X_5709_ _2414_ VPWR _2417_ VGND _2415_ _2416_ sg13g2_o21ai_1
XFILLER_3_804 VPWR VGND sg13g2_fill_1
XFILLER_12_66 VPWR VGND sg13g2_fill_2
Xhold171 mac2.products_ff\[146\] VPWR VGND net211 sg13g2_dlygate4sd3_1
Xhold160 mac2.sum_lvl1_ff\[9\] VPWR VGND net200 sg13g2_dlygate4sd3_1
Xhold193 mac2.sum_lvl2_ff\[42\] VPWR VGND net233 sg13g2_dlygate4sd3_1
Xhold182 mac2.sum_lvl1_ff\[79\] VPWR VGND net222 sg13g2_dlygate4sd3_1
XFILLER_37_85 VPWR VGND sg13g2_fill_2
XFILLER_15_911 VPWR VGND sg13g2_decap_4
XFILLER_42_752 VPWR VGND sg13g2_decap_4
XFILLER_15_966 VPWR VGND sg13g2_decap_8
XFILLER_30_969 VPWR VGND sg13g2_decap_8
X_4040_ _0844_ VPWR _0882_ VGND _0841_ _0845_ sg13g2_o21ai_1
X_5991_ net1043 VGND VPWR _0069_ mac1.products_ff\[0\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_17_281 VPWR VGND sg13g2_fill_2
XFILLER_33_730 VPWR VGND sg13g2_decap_8
X_4942_ _1743_ net850 net791 VPWR VGND sg13g2_nand2_1
X_4873_ _1681_ _1680_ _1652_ VPWR VGND sg13g2_nand2b_1
X_3824_ _0661_ _0669_ _0671_ _0672_ VPWR VGND sg13g2_or3_1
XFILLER_21_969 VPWR VGND sg13g2_decap_8
X_3755_ _0609_ net980 DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_6474_ net1012 VGND VPWR net453 mac2.total_sum\[2\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3686_ _0543_ net986 net1005 VPWR VGND sg13g2_nand2_1
X_5425_ mac1.sum_lvl3_ff\[33\] net341 _2186_ VPWR VGND sg13g2_and2_1
X_5356_ net480 _2132_ _0004_ VPWR VGND sg13g2_nor2b_2
X_5287_ VGND VPWR _2047_ _2069_ _2077_ _2071_ sg13g2_a21oi_1
X_4307_ _1131_ VPWR _1136_ VGND _1133_ _1134_ sg13g2_o21ai_1
X_4238_ _1066_ _1067_ _1061_ _1069_ VPWR VGND sg13g2_nand3_1
X_4169_ _0082_ _0988_ _1001_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_446 VPWR VGND sg13g2_fill_2
XFILLER_20_991 VPWR VGND sg13g2_decap_8
XFILLER_47_855 VPWR VGND sg13g2_decap_4
XFILLER_34_505 VPWR VGND sg13g2_decap_4
XFILLER_42_593 VPWR VGND sg13g2_decap_4
XFILLER_11_991 VPWR VGND sg13g2_decap_8
X_3540_ _0356_ _0399_ _0401_ VPWR VGND sg13g2_and2_1
X_3471_ _0331_ _0332_ _0326_ _0334_ VPWR VGND sg13g2_nand3_1
X_5210_ _2002_ _2003_ _2004_ VPWR VGND sg13g2_nor2b_1
X_6190_ net1082 VGND VPWR net49 mac1.sum_lvl2_ff\[11\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5141_ _1894_ _1891_ _1935_ _1937_ VPWR VGND sg13g2_a21o_1
X_5072_ _1869_ net789 net844 VPWR VGND sg13g2_nand2_1
X_4023_ _0866_ _0837_ _0864_ VPWR VGND sg13g2_xnor2_1
X_5974_ net808 _0256_ VPWR VGND sg13g2_buf_1
X_4925_ net799 net795 net851 net848 _1727_ VPWR VGND sg13g2_and4_1
X_4856_ VGND VPWR _1664_ _1665_ _1663_ _1604_ sg13g2_a21oi_2
X_3807_ _0647_ VPWR _0655_ VGND _0639_ _0649_ sg13g2_o21ai_1
XFILLER_21_799 VPWR VGND sg13g2_fill_1
X_4787_ _1596_ _1572_ _1598_ VPWR VGND sg13g2_xor2_1
X_3738_ _0593_ DP_2.matrix\[6\] net1011 VPWR VGND sg13g2_nand2_1
X_3669_ _0514_ _0526_ _0527_ VPWR VGND sg13g2_nor2_1
X_6457_ net1058 VGND VPWR net292 mac2.sum_lvl3_ff\[1\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_5408_ _2172_ mac1.sum_lvl3_ff\[30\] net377 VPWR VGND sg13g2_nand2_1
X_6388_ net1057 VGND VPWR net45 mac2.sum_lvl1_ff\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_5339_ _2118_ net538 _0001_ VPWR VGND sg13g2_xor2_1
XFILLER_28_343 VPWR VGND sg13g2_fill_2
XFILLER_29_888 VPWR VGND sg13g2_decap_8
XFILLER_43_324 VPWR VGND sg13g2_fill_1
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_11_243 VPWR VGND sg13g2_fill_1
XFILLER_4_954 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_58_clk clknet_4_9_0_clk clknet_leaf_58_clk VPWR VGND sg13g2_buf_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_15_560 VPWR VGND sg13g2_fill_2
X_5690_ _2396_ VPWR _2399_ VGND _2397_ _2398_ sg13g2_o21ai_1
XFILLER_30_541 VPWR VGND sg13g2_fill_1
X_4710_ _1521_ _1520_ _1486_ _1523_ VPWR VGND sg13g2_a21o_1
X_4641_ _1455_ _1449_ _1453_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_770 VPWR VGND sg13g2_fill_1
X_4572_ _1387_ _1369_ _0088_ VPWR VGND sg13g2_xor2_1
X_3523_ _0383_ _0382_ _0113_ VPWR VGND sg13g2_xor2_1
X_6311_ net1049 VGND VPWR net233 mac2.sum_lvl3_ff\[24\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_6242_ net1031 VGND VPWR net250 mac2.sum_lvl2_ff\[53\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3454_ _0317_ _0315_ _0316_ VPWR VGND sg13g2_nand2b_1
X_3385_ _2966_ _2963_ _2967_ VPWR VGND sg13g2_xor2_1
X_6173_ net1084 VGND VPWR net247 mac1.sum_lvl1_ff\[46\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5124_ _1920_ _1914_ _1919_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_49_clk clknet_4_10_0_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
X_5055_ _1813_ VPWR _1853_ VGND _1814_ _1815_ sg13g2_o21ai_1
X_4006_ _0847_ _0839_ _0849_ VPWR VGND sg13g2_xor2_1
XFILLER_38_674 VPWR VGND sg13g2_fill_1
XFILLER_38_1019 VPWR VGND sg13g2_decap_8
X_5957_ net865 _0231_ VPWR VGND sg13g2_buf_1
XFILLER_41_817 VPWR VGND sg13g2_decap_4
X_4908_ _1714_ _1701_ _1713_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_891 VPWR VGND sg13g2_decap_8
X_5888_ _2570_ VPWR _0226_ VGND net761 _2569_ sg13g2_o21ai_1
X_4839_ _1648_ _1642_ _1647_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_206 VPWR VGND sg13g2_fill_1
XFILLER_1_913 VPWR VGND sg13g2_decap_8
Xhold31 mac1.sum_lvl1_ff\[9\] VPWR VGND net71 sg13g2_dlygate4sd3_1
Xhold20 mac1.products_ff\[83\] VPWR VGND net60 sg13g2_dlygate4sd3_1
Xhold42 mac2.sum_lvl2_ff\[50\] VPWR VGND net82 sg13g2_dlygate4sd3_1
Xhold64 mac2.sum_lvl1_ff\[80\] VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold53 mac2.products_ff\[11\] VPWR VGND net93 sg13g2_dlygate4sd3_1
Xhold86 mac1.sum_lvl1_ff\[73\] VPWR VGND net126 sg13g2_dlygate4sd3_1
Xhold75 mac1.sum_lvl1_ff\[74\] VPWR VGND net115 sg13g2_dlygate4sd3_1
Xhold97 mac2.sum_lvl2_ff\[46\] VPWR VGND net137 sg13g2_dlygate4sd3_1
XFILLER_16_313 VPWR VGND sg13g2_fill_1
XFILLER_17_836 VPWR VGND sg13g2_fill_1
XFILLER_45_52 VPWR VGND sg13g2_fill_1
XFILLER_43_165 VPWR VGND sg13g2_fill_2
X_3170_ _2750_ VPWR _2762_ VGND _2758_ _2760_ sg13g2_o21ai_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_1017 VPWR VGND sg13g2_decap_8
Xfanout1040 net1042 net1040 VPWR VGND sg13g2_buf_8
XFILLER_0_990 VPWR VGND sg13g2_decap_8
Xfanout1062 net1063 net1062 VPWR VGND sg13g2_buf_8
Xfanout1051 net1053 net1051 VPWR VGND sg13g2_buf_8
Xfanout1073 net1074 net1073 VPWR VGND sg13g2_buf_8
XFILLER_48_961 VPWR VGND sg13g2_decap_8
Xfanout1095 net1097 net1095 VPWR VGND sg13g2_buf_8
Xfanout1084 net1087 net1084 VPWR VGND sg13g2_buf_8
XFILLER_47_493 VPWR VGND sg13g2_fill_2
X_5811_ _2517_ net784 net766 VPWR VGND sg13g2_nand2_1
XFILLER_16_880 VPWR VGND sg13g2_fill_2
XFILLER_35_699 VPWR VGND sg13g2_decap_8
X_5742_ DP_3.Q_range.out_data\[2\] DP_3.I_range.out_data\[2\] _2449_ VPWR VGND sg13g2_xor2_1
X_5673_ _2379_ VPWR _2382_ VGND _2380_ _2381_ sg13g2_o21ai_1
X_4624_ _1437_ _1436_ _1427_ _1439_ VPWR VGND sg13g2_a21o_1
Xhold501 _0061_ VPWR VGND net541 sg13g2_dlygate4sd3_1
X_4555_ _1356_ _1371_ _1372_ VPWR VGND sg13g2_nor2_1
X_3506_ _0368_ _0361_ _0366_ _0367_ VPWR VGND sg13g2_and3_1
X_4486_ _1310_ _1301_ _1309_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_1012 VPWR VGND sg13g2_decap_8
X_3437_ _0301_ _0294_ _0299_ _0300_ VPWR VGND sg13g2_and3_1
X_6225_ net1046 VGND VPWR net81 mac1.sum_lvl2_ff\[52\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6156_ net1054 VGND VPWR _0261_ DP_4.matrix\[73\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3368_ VGND VPWR _2936_ _2952_ _2953_ _2951_ sg13g2_a21oi_1
X_5107_ _1870_ VPWR _1903_ VGND _1867_ _1871_ sg13g2_o21ai_1
XFILLER_45_408 VPWR VGND sg13g2_fill_2
X_3299_ _2867_ VPWR _2887_ VGND _2864_ _2868_ sg13g2_o21ai_1
X_6087_ net1081 VGND VPWR _0211_ DP_2.matrix\[43\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_39_972 VPWR VGND sg13g2_decap_8
X_5038_ _1832_ _1833_ _1835_ _1836_ VPWR VGND sg13g2_or3_1
XFILLER_22_850 VPWR VGND sg13g2_fill_2
XFILLER_21_360 VPWR VGND sg13g2_fill_1
Xoutput32 net32 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_37_909 VPWR VGND sg13g2_decap_8
XFILLER_17_600 VPWR VGND sg13g2_fill_2
XFILLER_16_110 VPWR VGND sg13g2_fill_2
XFILLER_45_986 VPWR VGND sg13g2_decap_8
XFILLER_13_861 VPWR VGND sg13g2_fill_2
XFILLER_9_832 VPWR VGND sg13g2_fill_2
XFILLER_28_1007 VPWR VGND sg13g2_decap_8
X_4340_ _1168_ net870 net995 VPWR VGND sg13g2_nand2_1
X_4271_ _1096_ VPWR _1101_ VGND _1097_ _1099_ sg13g2_o21ai_1
X_6010_ net1067 VGND VPWR _0077_ mac1.products_ff\[71\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3222_ _2771_ _2768_ _2811_ _2813_ VPWR VGND sg13g2_a21o_1
X_3153_ _2745_ net892 net947 VPWR VGND sg13g2_nand2_1
XFILLER_28_909 VPWR VGND sg13g2_decap_8
X_3084_ _2678_ net944 net904 net946 net900 VPWR VGND sg13g2_a22oi_1
XFILLER_36_920 VPWR VGND sg13g2_decap_8
XFILLER_36_997 VPWR VGND sg13g2_decap_8
X_3986_ _0830_ _0797_ _0829_ VPWR VGND sg13g2_nand2b_1
X_5725_ net771 VPWR _2433_ VGND DP_2.matrix\[40\] net773 sg13g2_o21ai_1
X_5656_ _2364_ VPWR _2365_ VGND DP_1.I_range.out_data\[5\] _2359_ sg13g2_o21ai_1
X_4607_ _1422_ net885 net822 VPWR VGND sg13g2_nand2_1
X_5587_ _2310_ _2308_ net27 VPWR VGND sg13g2_xor2_1
Xhold320 mac2.sum_lvl2_ff\[3\] VPWR VGND net360 sg13g2_dlygate4sd3_1
Xhold331 DP_1.matrix\[38\] VPWR VGND net371 sg13g2_dlygate4sd3_1
Xhold353 mac1.sum_lvl3_ff\[11\] VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold342 _0049_ VPWR VGND net382 sg13g2_dlygate4sd3_1
X_4538_ _1356_ net886 net825 VPWR VGND sg13g2_nand2_1
Xhold364 DP_4.matrix\[5\] VPWR VGND net404 sg13g2_dlygate4sd3_1
Xfanout800 net282 net800 VPWR VGND sg13g2_buf_2
Xhold375 mac1.sum_lvl2_ff\[2\] VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold386 _0050_ VPWR VGND net426 sg13g2_dlygate4sd3_1
X_4469_ VGND VPWR _1234_ _1266_ _1294_ _1265_ sg13g2_a21oi_1
Xfanout822 net404 net822 VPWR VGND sg13g2_buf_8
X_6208_ net1083 VGND VPWR net242 mac1.sum_lvl2_ff\[32\] clknet_leaf_47_clk sg13g2_dfrbpq_2
Xhold397 _2270_ VPWR VGND net437 sg13g2_dlygate4sd3_1
Xfanout811 net331 net811 VPWR VGND sg13g2_buf_8
Xfanout833 net837 net833 VPWR VGND sg13g2_buf_8
Xfanout844 net845 net844 VPWR VGND sg13g2_buf_8
Xfanout855 net857 net855 VPWR VGND sg13g2_buf_2
Xfanout866 net473 net866 VPWR VGND sg13g2_buf_8
Xfanout877 DP_3.matrix\[5\] net877 VPWR VGND sg13g2_buf_8
XFILLER_46_717 VPWR VGND sg13g2_fill_2
Xfanout899 net902 net899 VPWR VGND sg13g2_buf_1
Xfanout888 net346 net888 VPWR VGND sg13g2_buf_1
X_6139_ net1096 VGND VPWR net76 mac1.sum_lvl1_ff\[14\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_27_931 VPWR VGND sg13g2_decap_8
XFILLER_14_603 VPWR VGND sg13g2_fill_1
XFILLER_42_945 VPWR VGND sg13g2_decap_8
XFILLER_14_669 VPWR VGND sg13g2_fill_1
XFILLER_41_444 VPWR VGND sg13g2_fill_1
XFILLER_9_128 VPWR VGND sg13g2_fill_2
XFILLER_42_31 VPWR VGND sg13g2_fill_1
XFILLER_37_706 VPWR VGND sg13g2_fill_2
XFILLER_18_997 VPWR VGND sg13g2_decap_8
XFILLER_33_923 VPWR VGND sg13g2_decap_8
X_3840_ _0670_ VPWR _0687_ VGND _0661_ _0671_ sg13g2_o21ai_1
X_3771_ _0620_ _0614_ _0076_ VPWR VGND sg13g2_xor2_1
X_5510_ mac2.sum_lvl3_ff\[21\] mac2.sum_lvl3_ff\[1\] _2251_ VPWR VGND sg13g2_nor2_1
XFILLER_9_673 VPWR VGND sg13g2_fill_1
X_6490_ net1026 VGND VPWR net7 DP_1.Q_range.out_data\[4\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5441_ _0039_ _2194_ _2197_ VPWR VGND sg13g2_xnor2_1
X_5372_ mac1.sum_lvl3_ff\[22\] mac1.sum_lvl3_ff\[2\] _2144_ VPWR VGND sg13g2_and2_1
XFILLER_5_890 VPWR VGND sg13g2_fill_1
X_4323_ VGND VPWR _1148_ _1149_ _1152_ _1130_ sg13g2_a21oi_1
X_4254_ _1084_ net870 net801 VPWR VGND sg13g2_nand2_1
X_3205_ _2796_ _2791_ _2795_ VPWR VGND sg13g2_xnor2_1
X_4185_ _1018_ _0998_ _1000_ VPWR VGND sg13g2_nand2_1
XFILLER_41_1004 VPWR VGND sg13g2_decap_8
X_3136_ _2728_ _2665_ _2729_ VPWR VGND sg13g2_xor2_1
X_3067_ _0094_ _2634_ _2661_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_967 VPWR VGND sg13g2_decap_8
X_5708_ net770 VPWR _2416_ VGND DP_2.matrix\[39\] net773 sg13g2_o21ai_1
X_3969_ VGND VPWR _0813_ _0812_ _0765_ sg13g2_or2_1
X_5639_ _2349_ _2350_ _2347_ _2352_ VPWR VGND sg13g2_nand3_1
Xhold161 mac1.sum_lvl1_ff\[78\] VPWR VGND net201 sg13g2_dlygate4sd3_1
Xhold150 mac2.sum_lvl1_ff\[78\] VPWR VGND net190 sg13g2_dlygate4sd3_1
Xhold172 mac1.products_ff\[140\] VPWR VGND net212 sg13g2_dlygate4sd3_1
Xhold194 mac2.products_ff\[139\] VPWR VGND net234 sg13g2_dlygate4sd3_1
Xhold183 mac2.products_ff\[2\] VPWR VGND net223 sg13g2_dlygate4sd3_1
XFILLER_46_547 VPWR VGND sg13g2_fill_2
XFILLER_2_1020 VPWR VGND sg13g2_decap_8
XFILLER_15_945 VPWR VGND sg13g2_decap_8
XFILLER_42_742 VPWR VGND sg13g2_fill_1
XFILLER_14_433 VPWR VGND sg13g2_fill_1
XFILLER_30_948 VPWR VGND sg13g2_decap_8
XFILLER_6_610 VPWR VGND sg13g2_decap_4
XFILLER_18_750 VPWR VGND sg13g2_fill_2
X_5990_ net1033 VGND VPWR net12 DP_3.Q_range.out_data\[6\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_4941_ _1728_ VPWR _1742_ VGND _1726_ _1729_ sg13g2_o21ai_1
X_4872_ _1678_ _1637_ _1680_ VPWR VGND sg13g2_xor2_1
X_3823_ VGND VPWR _0667_ _0668_ _0671_ _0662_ sg13g2_a21oi_1
XFILLER_21_948 VPWR VGND sg13g2_decap_8
X_3754_ _0595_ VPWR _0608_ VGND _0569_ _0593_ sg13g2_o21ai_1
X_6473_ net1013 VGND VPWR net475 mac2.total_sum\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3685_ _0511_ VPWR _0542_ VGND _0509_ _0512_ sg13g2_o21ai_1
X_5424_ VGND VPWR _2185_ net341 mac1.sum_lvl3_ff\[33\] sg13g2_or2_1
X_5355_ _2129_ net479 _2127_ _2132_ VPWR VGND sg13g2_nand3_1
X_5286_ _2073_ VPWR _2076_ VGND _2058_ _2075_ sg13g2_o21ai_1
X_4306_ _1131_ _1133_ _1134_ _1135_ VPWR VGND sg13g2_nor3_1
X_4237_ _1068_ _1061_ _1066_ _1067_ VPWR VGND sg13g2_and3_1
X_4168_ _0988_ _1001_ _1002_ VPWR VGND sg13g2_nor2b_1
X_3119_ _2712_ net941 net905 net944 net900 VPWR VGND sg13g2_a22oi_1
X_4099_ _0939_ _0938_ _0935_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_33 VPWR VGND sg13g2_fill_1
XFILLER_20_970 VPWR VGND sg13g2_decap_8
XFILLER_48_30 VPWR VGND sg13g2_fill_1
XFILLER_34_539 VPWR VGND sg13g2_fill_1
XFILLER_14_252 VPWR VGND sg13g2_fill_2
XFILLER_30_756 VPWR VGND sg13g2_decap_4
XFILLER_11_970 VPWR VGND sg13g2_decap_8
XFILLER_31_1025 VPWR VGND sg13g2_decap_4
XFILLER_10_491 VPWR VGND sg13g2_fill_1
XFILLER_7_985 VPWR VGND sg13g2_decap_8
X_3470_ _0333_ _0326_ _0331_ _0332_ VPWR VGND sg13g2_and3_1
XFILLER_43_4 VPWR VGND sg13g2_fill_2
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
X_5140_ VGND VPWR _1891_ _1894_ _1936_ _1935_ sg13g2_a21oi_1
X_5071_ _1868_ net787 net844 VPWR VGND sg13g2_nand2_1
X_4022_ _0865_ _0837_ _0864_ VPWR VGND sg13g2_nand2_1
X_5973_ net809 _0255_ VPWR VGND sg13g2_buf_1
X_4924_ _1726_ net852 net792 VPWR VGND sg13g2_nand2_1
XFILLER_20_233 VPWR VGND sg13g2_fill_2
X_4855_ _1632_ VPWR _1664_ VGND _1602_ _1631_ sg13g2_o21ai_1
X_3806_ _0653_ _0635_ _0078_ VPWR VGND sg13g2_xor2_1
X_4786_ _1597_ _1572_ _1596_ VPWR VGND sg13g2_nand2_1
X_3737_ _0592_ DP_2.matrix\[7\] net1010 VPWR VGND sg13g2_nand2_1
X_3668_ _0526_ _0516_ _0525_ VPWR VGND sg13g2_xnor2_1
X_6456_ net1058 VGND VPWR net268 mac2.sum_lvl3_ff\[0\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3599_ _0459_ _0443_ _0458_ VPWR VGND sg13g2_nand2_1
X_5407_ _2168_ VPWR _2171_ VGND _2167_ _2169_ sg13g2_o21ai_1
X_6387_ net1055 VGND VPWR net253 mac2.sum_lvl1_ff\[0\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_0_627 VPWR VGND sg13g2_decap_8
X_5338_ _2113_ _2117_ _2118_ VPWR VGND sg13g2_nor2_1
X_5269_ _2045_ _2037_ _2044_ _2060_ VPWR VGND sg13g2_a21o_1
XFILLER_29_867 VPWR VGND sg13g2_decap_8
XFILLER_31_509 VPWR VGND sg13g2_fill_1
XFILLER_11_222 VPWR VGND sg13g2_fill_2
XFILLER_4_933 VPWR VGND sg13g2_decap_8
XFILLER_38_119 VPWR VGND sg13g2_fill_1
XFILLER_47_642 VPWR VGND sg13g2_fill_1
XFILLER_35_859 VPWR VGND sg13g2_decap_8
XFILLER_15_572 VPWR VGND sg13g2_fill_1
XFILLER_43_892 VPWR VGND sg13g2_decap_8
XFILLER_30_531 VPWR VGND sg13g2_fill_1
X_4640_ _1449_ _1453_ _1454_ VPWR VGND sg13g2_and2_1
X_6310_ net1058 VGND VPWR net83 mac2.sum_lvl3_ff\[23\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4571_ _1369_ _1387_ _1388_ VPWR VGND sg13g2_and2_1
X_3522_ _0384_ _0382_ _0383_ VPWR VGND sg13g2_nand2_1
X_3453_ _0316_ DP_1.matrix\[0\] net926 VPWR VGND sg13g2_nand2_1
X_6241_ net1032 VGND VPWR net91 mac2.sum_lvl2_ff\[52\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_6172_ net1081 VGND VPWR net149 mac1.sum_lvl1_ff\[45\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_5123_ _1919_ _1868_ _1916_ VPWR VGND sg13g2_xnor2_1
X_3384_ _2964_ _2965_ _2966_ VPWR VGND sg13g2_nor2_1
XFILLER_29_119 VPWR VGND sg13g2_fill_1
X_5054_ _1851_ _1787_ _1852_ VPWR VGND sg13g2_xor2_1
X_4005_ _0847_ _0839_ _0848_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_314 VPWR VGND sg13g2_fill_1
XFILLER_37_152 VPWR VGND sg13g2_fill_2
XFILLER_26_859 VPWR VGND sg13g2_decap_8
XFILLER_34_870 VPWR VGND sg13g2_decap_8
X_5956_ net867 _0230_ VPWR VGND sg13g2_buf_1
X_4907_ _1713_ _1710_ _1712_ VPWR VGND sg13g2_xnor2_1
X_5887_ _2570_ net874 net761 VPWR VGND sg13g2_nand2_1
X_4838_ _1644_ _1646_ _1647_ VPWR VGND sg13g2_nor2_1
XFILLER_14_1020 VPWR VGND sg13g2_decap_8
X_4769_ _1579_ _1575_ _1580_ VPWR VGND sg13g2_xor2_1
XFILLER_4_229 VPWR VGND sg13g2_fill_1
X_6439_ net1093 VGND VPWR net124 mac2.sum_lvl2_ff\[15\] clknet_leaf_35_clk sg13g2_dfrbpq_1
XFILLER_20_56 VPWR VGND sg13g2_fill_1
XFILLER_1_969 VPWR VGND sg13g2_decap_8
XFILLER_0_457 VPWR VGND sg13g2_fill_2
Xhold21 mac1.products_ff\[8\] VPWR VGND net61 sg13g2_dlygate4sd3_1
Xhold32 mac2.sum_lvl1_ff\[41\] VPWR VGND net72 sg13g2_dlygate4sd3_1
Xhold10 mac2.sum_lvl1_ff\[10\] VPWR VGND net50 sg13g2_dlygate4sd3_1
Xhold54 mac1.sum_lvl1_ff\[12\] VPWR VGND net94 sg13g2_dlygate4sd3_1
Xhold43 mac2.sum_lvl2_ff\[41\] VPWR VGND net83 sg13g2_dlygate4sd3_1
XFILLER_29_631 VPWR VGND sg13g2_fill_1
Xhold65 mac2.sum_lvl1_ff\[7\] VPWR VGND net105 sg13g2_dlygate4sd3_1
Xhold87 mac1.sum_lvl1_ff\[7\] VPWR VGND net127 sg13g2_dlygate4sd3_1
Xhold76 mac1.sum_lvl1_ff\[39\] VPWR VGND net116 sg13g2_dlygate4sd3_1
Xhold98 mac2.products_ff\[69\] VPWR VGND net138 sg13g2_dlygate4sd3_1
XFILLER_28_152 VPWR VGND sg13g2_fill_1
XFILLER_16_336 VPWR VGND sg13g2_fill_1
XFILLER_17_859 VPWR VGND sg13g2_fill_2
XFILLER_45_86 VPWR VGND sg13g2_fill_1
XFILLER_12_553 VPWR VGND sg13g2_fill_1
XFILLER_12_575 VPWR VGND sg13g2_fill_1
XFILLER_4_763 VPWR VGND sg13g2_fill_1
Xfanout1030 net1038 net1030 VPWR VGND sg13g2_buf_8
XFILLER_48_940 VPWR VGND sg13g2_decap_8
Xfanout1074 net1075 net1074 VPWR VGND sg13g2_buf_8
Xfanout1041 net1042 net1041 VPWR VGND sg13g2_buf_8
Xfanout1063 net1098 net1063 VPWR VGND sg13g2_buf_8
Xfanout1052 net1053 net1052 VPWR VGND sg13g2_buf_8
Xfanout1085 net1086 net1085 VPWR VGND sg13g2_buf_8
Xfanout1096 net1097 net1096 VPWR VGND sg13g2_buf_8
XFILLER_47_472 VPWR VGND sg13g2_fill_1
XFILLER_35_612 VPWR VGND sg13g2_fill_1
XFILLER_35_645 VPWR VGND sg13g2_fill_2
X_5810_ _2516_ _2497_ _2515_ VPWR VGND sg13g2_nand2b_1
XFILLER_22_339 VPWR VGND sg13g2_fill_2
X_5741_ _2448_ DP_3.I_range.out_data\[2\] DP_3.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
X_5672_ net772 VPWR _2381_ VGND net972 net774 sg13g2_o21ai_1
X_4623_ _1436_ _1437_ _1427_ _1438_ VPWR VGND sg13g2_nand3_1
Xhold502 mac2.sum_lvl2_ff\[9\] VPWR VGND net542 sg13g2_dlygate4sd3_1
X_4554_ _1371_ net885 net824 VPWR VGND sg13g2_nand2_1
X_3505_ _0362_ VPWR _0367_ VGND _0363_ _0365_ sg13g2_o21ai_1
X_4485_ _1309_ _1272_ _1307_ VPWR VGND sg13g2_xnor2_1
X_6224_ net1049 VGND VPWR net170 mac1.sum_lvl2_ff\[51\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3436_ _0295_ VPWR _0300_ VGND _0296_ _0298_ sg13g2_o21ai_1
X_6155_ net1054 VGND VPWR _0260_ DP_4.matrix\[72\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3367_ _2952_ _2936_ _0099_ VPWR VGND sg13g2_xor2_1
X_6086_ net1081 VGND VPWR _0210_ DP_2.matrix\[42\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5106_ _1861_ VPWR _1902_ VGND _1819_ _1859_ sg13g2_o21ai_1
X_5037_ _1835_ net839 net797 net842 net793 VPWR VGND sg13g2_a22oi_1
X_3298_ _2886_ _2885_ _2883_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_951 VPWR VGND sg13g2_decap_8
XFILLER_38_472 VPWR VGND sg13g2_decap_8
XFILLER_25_100 VPWR VGND sg13g2_fill_2
X_5939_ net920 _0205_ VPWR VGND sg13g2_buf_1
XFILLER_22_862 VPWR VGND sg13g2_fill_1
XFILLER_40_158 VPWR VGND sg13g2_decap_8
XFILLER_40_169 VPWR VGND sg13g2_fill_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_210 VPWR VGND sg13g2_fill_2
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_0_276 VPWR VGND sg13g2_fill_1
XFILLER_45_965 VPWR VGND sg13g2_decap_8
XFILLER_29_494 VPWR VGND sg13g2_decap_4
XFILLER_13_840 VPWR VGND sg13g2_fill_1
XFILLER_31_147 VPWR VGND sg13g2_fill_2
X_4270_ _1096_ _1097_ _1099_ _1100_ VPWR VGND sg13g2_or3_1
X_3221_ VGND VPWR _2768_ _2771_ _2812_ _2811_ sg13g2_a21oi_1
X_3152_ _2744_ net953 net890 VPWR VGND sg13g2_nand2_1
X_3083_ net900 net946 net904 _2677_ VPWR VGND net944 sg13g2_nand4_1
XFILLER_35_453 VPWR VGND sg13g2_fill_2
XFILLER_36_976 VPWR VGND sg13g2_decap_8
X_3985_ _0829_ _0798_ _0827_ VPWR VGND sg13g2_xnor2_1
X_5724_ net928 net775 _2432_ VPWR VGND sg13g2_nor2_1
X_5655_ DP_1.I_range.out_data\[6\] DP_1.I_range.out_data\[4\] DP_1.Q_range.out_data\[4\]
+ _2363_ _2364_ VPWR VGND sg13g2_nor4_1
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
X_4606_ _1404_ VPWR _1421_ VGND _1395_ _1405_ sg13g2_o21ai_1
Xhold310 DP_4.matrix\[3\] VPWR VGND net350 sg13g2_dlygate4sd3_1
X_5586_ mac2.total_sum\[2\] mac1.total_sum\[2\] _2310_ VPWR VGND sg13g2_xor2_1
Xhold343 mac1.sum_lvl3_ff\[3\] VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold321 _2203_ VPWR VGND net361 sg13g2_dlygate4sd3_1
X_4537_ _1354_ _1348_ _0086_ VPWR VGND sg13g2_xor2_1
Xhold332 DP_3.matrix\[73\] VPWR VGND net372 sg13g2_dlygate4sd3_1
Xhold387 DP_2.matrix\[0\] VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold376 _2090_ VPWR VGND net416 sg13g2_dlygate4sd3_1
Xhold365 mac1.sum_lvl3_ff\[8\] VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold354 _2176_ VPWR VGND net394 sg13g2_dlygate4sd3_1
X_4468_ _1291_ _1290_ _1293_ VPWR VGND sg13g2_xor2_1
Xfanout801 net802 net801 VPWR VGND sg13g2_buf_8
Xfanout823 net824 net823 VPWR VGND sg13g2_buf_8
X_3419_ _0284_ _0282_ _0283_ VPWR VGND sg13g2_nand2_1
X_6207_ net1083 VGND VPWR net220 mac1.sum_lvl2_ff\[31\] clknet_leaf_47_clk sg13g2_dfrbpq_2
Xhold398 _2276_ VPWR VGND net438 sg13g2_dlygate4sd3_1
Xfanout812 DP_4.matrix\[38\] net812 VPWR VGND sg13g2_buf_1
Xfanout834 net837 net834 VPWR VGND sg13g2_buf_1
Xfanout856 net857 net856 VPWR VGND sg13g2_buf_8
Xfanout867 net327 net867 VPWR VGND sg13g2_buf_8
X_6138_ net1060 VGND VPWR _0245_ DP_4.matrix\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_4399_ _1226_ _1218_ _1225_ VPWR VGND sg13g2_xnor2_1
Xfanout845 DP_3.matrix\[77\] net845 VPWR VGND sg13g2_buf_8
XFILLER_46_707 VPWR VGND sg13g2_fill_1
Xfanout889 DP_2.matrix\[78\] net889 VPWR VGND sg13g2_buf_8
Xfanout878 net879 net878 VPWR VGND sg13g2_buf_8
X_6069_ net1045 VGND VPWR _0199_ DP_2.matrix\[3\] clknet_leaf_56_clk sg13g2_dfrbpq_2
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_42_924 VPWR VGND sg13g2_decap_8
XFILLER_13_169 VPWR VGND sg13g2_fill_2
XFILLER_42_43 VPWR VGND sg13g2_decap_4
XFILLER_10_865 VPWR VGND sg13g2_fill_2
XFILLER_6_847 VPWR VGND sg13g2_fill_1
XFILLER_10_898 VPWR VGND sg13g2_fill_1
XFILLER_49_567 VPWR VGND sg13g2_fill_1
XFILLER_18_976 VPWR VGND sg13g2_decap_8
XFILLER_33_902 VPWR VGND sg13g2_decap_8
XFILLER_45_784 VPWR VGND sg13g2_fill_2
XFILLER_33_979 VPWR VGND sg13g2_decap_8
X_3770_ _0621_ _0614_ _0620_ VPWR VGND sg13g2_nand2_1
XFILLER_32_467 VPWR VGND sg13g2_decap_8
XFILLER_41_990 VPWR VGND sg13g2_decap_8
XFILLER_12_191 VPWR VGND sg13g2_fill_1
X_5440_ mac2.sum_lvl2_ff\[1\] mac2.sum_lvl2_ff\[20\] _2197_ VPWR VGND sg13g2_xor2_1
X_5371_ _2140_ VPWR _2143_ VGND _2139_ _2141_ sg13g2_o21ai_1
XFILLER_5_880 VPWR VGND sg13g2_fill_1
X_4322_ _1148_ _1149_ _1130_ _1151_ VPWR VGND sg13g2_nand3_1
X_4253_ _1083_ net801 DP_3.matrix\[36\] net803 net869 VPWR VGND sg13g2_a22oi_1
X_3204_ _2795_ _2745_ _2792_ VPWR VGND sg13g2_xnor2_1
X_4184_ _1016_ _1006_ _1017_ VPWR VGND sg13g2_xor2_1
X_3135_ _2728_ _2725_ _2727_ VPWR VGND sg13g2_nand2_1
X_3066_ _2661_ _2660_ _2659_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_423 VPWR VGND sg13g2_fill_2
XFILLER_24_946 VPWR VGND sg13g2_decap_8
XFILLER_35_261 VPWR VGND sg13g2_fill_2
XFILLER_23_434 VPWR VGND sg13g2_fill_2
X_3968_ _0812_ net914 net963 VPWR VGND sg13g2_nand2_1
X_5707_ net929 net775 _2415_ VPWR VGND sg13g2_nor2_1
XFILLER_32_990 VPWR VGND sg13g2_decap_8
X_3899_ _0743_ _0744_ _0714_ _0745_ VPWR VGND sg13g2_nand3_1
X_5638_ VGND VPWR _2347_ _2349_ _2351_ _2350_ sg13g2_a21oi_1
XFILLER_3_817 VPWR VGND sg13g2_decap_8
X_5569_ net400 _2297_ _0052_ VPWR VGND sg13g2_nor2b_1
Xhold162 mac1.products_ff\[148\] VPWR VGND net202 sg13g2_dlygate4sd3_1
Xhold140 mac1.sum_lvl1_ff\[81\] VPWR VGND net180 sg13g2_dlygate4sd3_1
Xhold151 mac2.products_ff\[78\] VPWR VGND net191 sg13g2_dlygate4sd3_1
Xhold184 mac1.products_ff\[68\] VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold173 mac1.sum_lvl1_ff\[87\] VPWR VGND net213 sg13g2_dlygate4sd3_1
Xhold195 mac2.sum_lvl1_ff\[73\] VPWR VGND net235 sg13g2_dlygate4sd3_1
XFILLER_18_239 VPWR VGND sg13g2_fill_2
XFILLER_18_1018 VPWR VGND sg13g2_decap_8
XFILLER_30_927 VPWR VGND sg13g2_decap_8
XFILLER_49_342 VPWR VGND sg13g2_fill_2
XFILLER_49_331 VPWR VGND sg13g2_fill_2
XFILLER_49_386 VPWR VGND sg13g2_fill_1
X_4940_ VGND VPWR _1741_ _1740_ _1738_ sg13g2_or2_1
X_4871_ _1637_ _1678_ _1679_ VPWR VGND sg13g2_nor2_1
XFILLER_45_592 VPWR VGND sg13g2_decap_4
XFILLER_17_283 VPWR VGND sg13g2_fill_1
X_3822_ _0667_ _0668_ _0662_ _0670_ VPWR VGND sg13g2_nand3_1
XFILLER_21_927 VPWR VGND sg13g2_decap_8
XFILLER_33_787 VPWR VGND sg13g2_fill_1
X_3753_ VGND VPWR _0577_ _0599_ _0607_ _0601_ sg13g2_a21oi_1
X_6472_ net1012 VGND VPWR net306 mac2.total_sum\[0\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3684_ _0522_ VPWR _0541_ VGND _0476_ _0520_ sg13g2_o21ai_1
X_5423_ _2181_ VPWR _2184_ VGND _2180_ _2182_ sg13g2_o21ai_1
X_5354_ VGND VPWR _2127_ _2129_ _2131_ net479 sg13g2_a21oi_1
X_4305_ _1134_ net861 net809 net808 net864 VPWR VGND sg13g2_a22oi_1
X_5285_ _0154_ _2058_ _2074_ VPWR VGND sg13g2_xnor2_1
X_4236_ _1062_ VPWR _1067_ VGND _1063_ _1065_ sg13g2_o21ai_1
X_4167_ _1001_ _0989_ _0999_ VPWR VGND sg13g2_xnor2_1
X_3118_ net900 net944 net905 _2711_ VPWR VGND net941 sg13g2_nand4_1
X_4098_ _0937_ _0909_ _0938_ VPWR VGND sg13g2_xor2_1
X_3049_ net905 net899 net949 net946 _2644_ VPWR VGND sg13g2_and4_1
XFILLER_11_448 VPWR VGND sg13g2_fill_1
XFILLER_19_504 VPWR VGND sg13g2_fill_2
XFILLER_42_540 VPWR VGND sg13g2_fill_2
XFILLER_31_1004 VPWR VGND sg13g2_decap_8
XFILLER_7_964 VPWR VGND sg13g2_decap_8
X_5070_ _1867_ net848 net785 VPWR VGND sg13g2_nand2_1
XFILLER_49_150 VPWR VGND sg13g2_fill_2
X_4021_ _0862_ _0838_ _0864_ VPWR VGND sg13g2_xor2_1
XFILLER_37_356 VPWR VGND sg13g2_fill_2
XFILLER_38_879 VPWR VGND sg13g2_decap_8
X_5972_ net811 _0254_ VPWR VGND sg13g2_buf_1
XFILLER_18_581 VPWR VGND sg13g2_fill_2
X_4923_ VGND VPWR _1718_ _1721_ _1725_ _1719_ sg13g2_a21oi_1
XFILLER_33_573 VPWR VGND sg13g2_fill_1
X_4854_ _1605_ _1662_ _1663_ VPWR VGND sg13g2_nor2b_1
X_3805_ _0635_ _0653_ _0654_ VPWR VGND sg13g2_and2_1
X_4785_ _1595_ _1583_ _1596_ VPWR VGND sg13g2_xor2_1
X_3736_ _0591_ net982 net1005 VPWR VGND sg13g2_nand2_1
X_6455_ net1096 VGND VPWR net63 mac2.sum_lvl2_ff\[34\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3667_ _0525_ _0517_ _0523_ VPWR VGND sg13g2_xnor2_1
X_6386_ net1032 VGND VPWR _0155_ mac2.products_ff\[151\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5406_ _0031_ _2167_ net294 VPWR VGND sg13g2_xnor2_1
X_3598_ _0457_ _0450_ _0458_ VPWR VGND sg13g2_xor2_1
X_5337_ VPWR VGND mac1.sum_lvl2_ff\[9\] _2110_ mac1.sum_lvl2_ff\[28\] mac1.sum_lvl2_ff\[27\]
+ _2117_ mac1.sum_lvl2_ff\[8\] sg13g2_a221oi_1
X_5268_ _2049_ _2051_ _2059_ VPWR VGND sg13g2_and2_1
X_4219_ _1027_ VPWR _1050_ VGND _1004_ _1025_ sg13g2_o21ai_1
X_5199_ _1993_ _1988_ _1991_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_345 VPWR VGND sg13g2_fill_1
XFILLER_24_595 VPWR VGND sg13g2_decap_4
XFILLER_11_267 VPWR VGND sg13g2_fill_2
XFILLER_4_989 VPWR VGND sg13g2_decap_8
XFILLER_47_610 VPWR VGND sg13g2_fill_1
XFILLER_19_312 VPWR VGND sg13g2_fill_1
XFILLER_43_871 VPWR VGND sg13g2_decap_8
XFILLER_15_562 VPWR VGND sg13g2_fill_1
X_4570_ _1385_ _1384_ _1387_ VPWR VGND sg13g2_xor2_1
X_3521_ _0343_ VPWR _0383_ VGND _0344_ _0345_ sg13g2_o21ai_1
X_3452_ _0292_ VPWR _0315_ VGND _0269_ _0290_ sg13g2_o21ai_1
X_6240_ net1034 VGND VPWR net243 mac2.sum_lvl2_ff\[51\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3383_ _2965_ net989 net940 net936 net991 VPWR VGND sg13g2_a22oi_1
X_6171_ net1080 VGND VPWR net240 mac1.sum_lvl1_ff\[44\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5122_ _1868_ _1916_ _1918_ VPWR VGND sg13g2_and2_1
X_5053_ _1851_ _1848_ _1850_ VPWR VGND sg13g2_nand2_1
X_4004_ _0847_ _0840_ _0846_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_827 VPWR VGND sg13g2_fill_2
XFILLER_26_838 VPWR VGND sg13g2_decap_8
X_5955_ net869 _0229_ VPWR VGND sg13g2_buf_1
X_4906_ _1712_ _1695_ _1711_ VPWR VGND sg13g2_xnor2_1
X_5886_ _2482_ _2478_ _2569_ VPWR VGND sg13g2_xor2_1
X_4837_ _1646_ DP_4.matrix\[7\] net877 net821 net875 VPWR VGND sg13g2_a22oi_1
XFILLER_21_598 VPWR VGND sg13g2_fill_1
X_4768_ _1579_ _1536_ _1577_ VPWR VGND sg13g2_xnor2_1
X_3719_ _0575_ _0539_ _0573_ VPWR VGND sg13g2_xnor2_1
X_4699_ _1512_ _1505_ _1510_ _1511_ VPWR VGND sg13g2_and3_1
X_6438_ net1093 VGND VPWR net178 mac2.sum_lvl2_ff\[14\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_6369_ net1094 VGND VPWR _0132_ mac2.products_ff\[82\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_1_948 VPWR VGND sg13g2_decap_8
XFILLER_49_919 VPWR VGND sg13g2_decap_8
Xhold11 mac1.products_ff\[137\] VPWR VGND net51 sg13g2_dlygate4sd3_1
Xhold22 mac2.products_ff\[77\] VPWR VGND net62 sg13g2_dlygate4sd3_1
Xhold44 mac2.sum_lvl1_ff\[75\] VPWR VGND net84 sg13g2_dlygate4sd3_1
XFILLER_29_610 VPWR VGND sg13g2_fill_2
Xhold55 mac2.sum_lvl1_ff\[76\] VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold33 mac2.sum_lvl1_ff\[46\] VPWR VGND net73 sg13g2_dlygate4sd3_1
Xhold66 mac1.sum_lvl2_ff\[44\] VPWR VGND net106 sg13g2_dlygate4sd3_1
XFILLER_21_1025 VPWR VGND sg13g2_decap_4
Xhold77 mac2.sum_lvl2_ff\[44\] VPWR VGND net117 sg13g2_dlygate4sd3_1
Xhold99 mac2.sum_lvl1_ff\[36\] VPWR VGND net139 sg13g2_dlygate4sd3_1
Xhold88 mac2.sum_lvl1_ff\[84\] VPWR VGND net128 sg13g2_dlygate4sd3_1
XFILLER_40_885 VPWR VGND sg13g2_decap_8
XFILLER_8_558 VPWR VGND sg13g2_fill_1
Xfanout1031 net1034 net1031 VPWR VGND sg13g2_buf_8
Xfanout1020 net1021 net1020 VPWR VGND sg13g2_buf_8
Xfanout1064 net1066 net1064 VPWR VGND sg13g2_buf_8
Xfanout1042 net1063 net1042 VPWR VGND sg13g2_buf_8
Xfanout1053 net1063 net1053 VPWR VGND sg13g2_buf_8
Xfanout1086 net1087 net1086 VPWR VGND sg13g2_buf_8
Xfanout1097 net1098 net1097 VPWR VGND sg13g2_buf_8
Xfanout1075 net1077 net1075 VPWR VGND sg13g2_buf_8
XFILLER_48_996 VPWR VGND sg13g2_decap_8
XFILLER_19_197 VPWR VGND sg13g2_fill_2
X_5740_ _2447_ _2445_ _2446_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_1021 VPWR VGND sg13g2_decap_8
XFILLER_31_852 VPWR VGND sg13g2_fill_2
X_5671_ net987 net776 _2380_ VPWR VGND sg13g2_nor2_1
XFILLER_30_373 VPWR VGND sg13g2_fill_2
XFILLER_31_885 VPWR VGND sg13g2_decap_8
X_4622_ _1434_ _1433_ _1428_ _1437_ VPWR VGND sg13g2_a21o_1
X_4553_ _1370_ net824 net886 net825 net884 VPWR VGND sg13g2_a22oi_1
X_4484_ _1272_ _1307_ _1308_ VPWR VGND sg13g2_nor2b_1
X_3504_ _0362_ _0363_ _0365_ _0366_ VPWR VGND sg13g2_or3_1
Xhold503 _2224_ VPWR VGND net543 sg13g2_dlygate4sd3_1
X_3435_ _0295_ _0296_ _0298_ _0299_ VPWR VGND sg13g2_or3_1
X_6223_ net1024 VGND VPWR net236 mac1.sum_lvl2_ff\[50\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_6154_ net1095 VGND VPWR _0259_ DP_4.matrix\[43\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3366_ _2950_ _2937_ _2952_ VPWR VGND sg13g2_xor2_1
X_3297_ VGND VPWR _2885_ _2884_ _2833_ sg13g2_or2_1
X_6085_ net1021 VGND VPWR _0097_ mac1.products_ff\[148\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5105_ _1887_ VPWR _1901_ VGND _1865_ _1888_ sg13g2_o21ai_1
XFILLER_39_930 VPWR VGND sg13g2_decap_8
X_5036_ net793 net842 net797 _1834_ VPWR VGND net839 sg13g2_nand4_1
X_5938_ net923 _0204_ VPWR VGND sg13g2_buf_1
XFILLER_41_627 VPWR VGND sg13g2_fill_2
XFILLER_22_852 VPWR VGND sg13g2_fill_1
X_5869_ _2557_ VPWR _0203_ VGND _2443_ _2558_ sg13g2_o21ai_1
Xoutput23 net23 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_233 VPWR VGND sg13g2_fill_1
XFILLER_17_602 VPWR VGND sg13g2_fill_1
XFILLER_45_944 VPWR VGND sg13g2_decap_8
XFILLER_16_112 VPWR VGND sg13g2_fill_1
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_13_863 VPWR VGND sg13g2_fill_1
X_3220_ _2809_ _2777_ _2811_ VPWR VGND sg13g2_xor2_1
X_3151_ _2716_ VPWR _2743_ VGND _2707_ _2717_ sg13g2_o21ai_1
XFILLER_48_771 VPWR VGND sg13g2_decap_8
X_3082_ net904 net901 net946 net944 _2676_ VPWR VGND sg13g2_and4_1
XFILLER_35_410 VPWR VGND sg13g2_fill_1
XFILLER_36_955 VPWR VGND sg13g2_decap_8
XFILLER_23_616 VPWR VGND sg13g2_decap_4
X_3984_ _0828_ _0798_ _0827_ VPWR VGND sg13g2_nand2_1
X_5723_ _2431_ net893 net763 VPWR VGND sg13g2_nand2_1
X_5654_ DP_1.Q_range.out_data\[3\] _2362_ _2363_ VPWR VGND DP_1.I_range.out_data\[3\]
+ sg13g2_nand3b_1
X_4605_ _1418_ _1417_ _1420_ VPWR VGND sg13g2_xor2_1
X_5585_ mac1.total_sum\[2\] mac2.total_sum\[2\] _2309_ VPWR VGND sg13g2_and2_1
Xhold300 _0063_ VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold311 _0247_ VPWR VGND net351 sg13g2_dlygate4sd3_1
Xhold344 _2148_ VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold333 mac1.sum_lvl3_ff\[14\] VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold322 _0041_ VPWR VGND net362 sg13g2_dlygate4sd3_1
X_4536_ _1355_ _1348_ _1354_ VPWR VGND sg13g2_nand2_1
X_4467_ VGND VPWR _1292_ _1291_ _1290_ sg13g2_or2_1
Xhold366 _2164_ VPWR VGND net406 sg13g2_dlygate4sd3_1
Xhold377 _0008_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold355 _0018_ VPWR VGND net395 sg13g2_dlygate4sd3_1
Xfanout802 net465 net802 VPWR VGND sg13g2_buf_8
Xfanout824 net344 net824 VPWR VGND sg13g2_buf_8
Xhold388 DP_4.matrix\[7\] VPWR VGND net428 sg13g2_dlygate4sd3_1
X_4398_ _1223_ _1224_ _1225_ VPWR VGND sg13g2_nor2b_1
X_3418_ _0283_ _2978_ _2980_ VPWR VGND sg13g2_nand2_1
X_6206_ net1084 VGND VPWR net221 mac1.sum_lvl2_ff\[30\] clknet_leaf_48_clk sg13g2_dfrbpq_1
Xhold399 _0062_ VPWR VGND net439 sg13g2_dlygate4sd3_1
Xfanout813 net330 net813 VPWR VGND sg13g2_buf_8
Xfanout857 net447 net857 VPWR VGND sg13g2_buf_8
X_3349_ VGND VPWR _2905_ _2930_ _2935_ _2931_ sg13g2_a21oi_1
X_6137_ net1055 VGND VPWR _0244_ DP_4.matrix\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_1
Xfanout835 net837 net835 VPWR VGND sg13g2_buf_2
Xfanout846 net847 net846 VPWR VGND sg13g2_buf_8
Xfanout879 net517 net879 VPWR VGND sg13g2_buf_8
Xfanout868 DP_3.matrix\[38\] net868 VPWR VGND sg13g2_buf_2
XFILLER_46_719 VPWR VGND sg13g2_fill_1
X_6068_ net1046 VGND VPWR net389 DP_2.matrix\[2\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5019_ _1794_ VPWR _1817_ VGND _1759_ _1792_ sg13g2_o21ai_1
XFILLER_42_903 VPWR VGND sg13g2_decap_8
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_14_616 VPWR VGND sg13g2_fill_2
XFILLER_26_476 VPWR VGND sg13g2_fill_2
XFILLER_41_457 VPWR VGND sg13g2_fill_1
XFILLER_42_99 VPWR VGND sg13g2_decap_4
XFILLER_5_369 VPWR VGND sg13g2_fill_2
XFILLER_1_520 VPWR VGND sg13g2_fill_2
XFILLER_49_546 VPWR VGND sg13g2_decap_8
XFILLER_49_579 VPWR VGND sg13g2_decap_8
XFILLER_36_207 VPWR VGND sg13g2_fill_2
XFILLER_37_708 VPWR VGND sg13g2_fill_1
XFILLER_18_955 VPWR VGND sg13g2_decap_8
XFILLER_33_958 VPWR VGND sg13g2_decap_8
XFILLER_34_1024 VPWR VGND sg13g2_decap_4
XFILLER_9_642 VPWR VGND sg13g2_fill_2
XFILLER_9_631 VPWR VGND sg13g2_fill_1
X_5370_ _0023_ _2139_ _2142_ VPWR VGND sg13g2_xnor2_1
X_4321_ _1150_ _1130_ _1148_ _1149_ VPWR VGND sg13g2_and3_1
X_4252_ _1059_ VPWR _1082_ VGND _1024_ _1057_ sg13g2_o21ai_1
X_3203_ _2745_ _2792_ _2794_ VPWR VGND sg13g2_and2_1
X_4183_ _1016_ _1014_ _1015_ VPWR VGND sg13g2_nand2_1
X_3134_ _2724_ _2723_ _2694_ _2727_ VPWR VGND sg13g2_a21o_1
X_3065_ _2632_ VPWR _2660_ VGND _2656_ _2657_ sg13g2_o21ai_1
XFILLER_36_741 VPWR VGND sg13g2_decap_4
X_3967_ _0811_ net968 net910 VPWR VGND sg13g2_nand2_1
X_5706_ _2414_ net895 net763 VPWR VGND sg13g2_nand2_1
X_3898_ _0721_ VPWR _0744_ VGND _0740_ _0742_ sg13g2_o21ai_1
Xclkbuf_leaf_30_clk clknet_4_12_0_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_5637_ _2350_ mac1.total_sum\[13\] mac2.total_sum\[13\] VPWR VGND sg13g2_xnor2_1
X_5568_ _2294_ net399 _2292_ _2297_ VPWR VGND sg13g2_nand3_1
X_4519_ VGND VPWR _1311_ _1334_ _1341_ _1336_ sg13g2_a21oi_1
Xhold141 mac1.sum_lvl2_ff\[38\] VPWR VGND net181 sg13g2_dlygate4sd3_1
Xhold152 mac1.sum_lvl1_ff\[44\] VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold130 mac1.sum_lvl1_ff\[85\] VPWR VGND net170 sg13g2_dlygate4sd3_1
Xhold185 mac1.products_ff\[146\] VPWR VGND net225 sg13g2_dlygate4sd3_1
Xhold163 mac2.products_ff\[70\] VPWR VGND net203 sg13g2_dlygate4sd3_1
Xhold174 mac2.products_ff\[72\] VPWR VGND net214 sg13g2_dlygate4sd3_1
X_5499_ VGND VPWR mac2.sum_lvl2_ff\[32\] mac2.sum_lvl2_ff\[13\] _2243_ _2241_ sg13g2_a21oi_1
Xhold196 mac1.sum_lvl1_ff\[84\] VPWR VGND net236 sg13g2_dlygate4sd3_1
XFILLER_46_538 VPWR VGND sg13g2_fill_2
XFILLER_42_711 VPWR VGND sg13g2_fill_1
XFILLER_30_906 VPWR VGND sg13g2_decap_8
XFILLER_23_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_4_5_0_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_5_122 VPWR VGND sg13g2_fill_1
XFILLER_5_144 VPWR VGND sg13g2_fill_2
XFILLER_18_752 VPWR VGND sg13g2_fill_1
X_4870_ _1678_ _1669_ _1677_ VPWR VGND sg13g2_xnor2_1
X_3821_ _0669_ _0662_ _0667_ _0668_ VPWR VGND sg13g2_and3_1
X_3752_ _0603_ VPWR _0606_ VGND _0588_ _0605_ sg13g2_o21ai_1
Xclkbuf_leaf_12_clk clknet_4_6_0_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_6471_ net1037 VGND VPWR _0038_ mac2.sum_lvl3_ff\[15\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3683_ _0540_ _0539_ _0537_ VPWR VGND sg13g2_nand2b_1
X_5422_ _0019_ _2180_ net324 VPWR VGND sg13g2_xnor2_1
X_5353_ _2130_ mac1.sum_lvl2_ff\[32\] net478 VPWR VGND sg13g2_xnor2_1
X_4304_ net809 DP_3.matrix\[40\] net807 DP_3.matrix\[41\] _1133_ VPWR VGND sg13g2_and4_1
X_5284_ VPWR _2075_ _2074_ VGND sg13g2_inv_1
X_4235_ _1062_ _1063_ _1065_ _1066_ VPWR VGND sg13g2_or3_1
X_4166_ _1000_ _0999_ _0989_ VPWR VGND sg13g2_nand2b_1
X_3117_ net905 net900 net944 net941 _2710_ VPWR VGND sg13g2_and4_1
XFILLER_28_549 VPWR VGND sg13g2_fill_2
XFILLER_43_508 VPWR VGND sg13g2_fill_2
X_4097_ _0937_ net909 net962 VPWR VGND sg13g2_nand2_1
X_3048_ _2643_ net896 net952 VPWR VGND sg13g2_nand2_1
XFILLER_36_582 VPWR VGND sg13g2_fill_2
XFILLER_23_243 VPWR VGND sg13g2_fill_1
XFILLER_11_416 VPWR VGND sg13g2_fill_2
X_4999_ net797 net793 net844 net841 _1798_ VPWR VGND sg13g2_and4_1
XFILLER_3_648 VPWR VGND sg13g2_fill_2
XFILLER_24_1023 VPWR VGND sg13g2_decap_4
XFILLER_47_869 VPWR VGND sg13g2_decap_8
XFILLER_46_368 VPWR VGND sg13g2_fill_2
XFILLER_15_700 VPWR VGND sg13g2_fill_1
XFILLER_15_733 VPWR VGND sg13g2_fill_1
XFILLER_7_910 VPWR VGND sg13g2_fill_2
XFILLER_7_943 VPWR VGND sg13g2_decap_8
XFILLER_43_6 VPWR VGND sg13g2_fill_1
XFILLER_49_140 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_1_191 VPWR VGND sg13g2_fill_1
X_4020_ _0863_ _0838_ _0862_ VPWR VGND sg13g2_nand2_1
XFILLER_25_519 VPWR VGND sg13g2_decap_8
X_5971_ net813 _0253_ VPWR VGND sg13g2_buf_1
X_4922_ _1724_ net854 net790 VPWR VGND sg13g2_nand2_1
X_4853_ VGND VPWR _1601_ _1632_ _1662_ _1631_ sg13g2_a21oi_1
X_4784_ _1593_ _1584_ _1595_ VPWR VGND sg13g2_xor2_1
X_3804_ _0651_ _0650_ _0653_ VPWR VGND sg13g2_xor2_1
X_3735_ _0575_ _0567_ _0574_ _0590_ VPWR VGND sg13g2_a21o_1
X_6454_ net1097 VGND VPWR net118 mac2.sum_lvl2_ff\[33\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_5405_ net293 mac1.sum_lvl3_ff\[29\] _2170_ VPWR VGND sg13g2_xor2_1
X_3666_ _0524_ _0517_ _0523_ VPWR VGND sg13g2_nand2_1
X_6385_ net1031 VGND VPWR _0154_ mac2.products_ff\[150\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3597_ _0457_ _0451_ _0455_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_1023 VPWR VGND sg13g2_decap_4
X_5336_ net537 mac1.sum_lvl2_ff\[29\] _2116_ VPWR VGND sg13g2_xor2_1
X_5267_ VPWR VGND _2034_ _2053_ _2057_ _2029_ _2058_ _2054_ sg13g2_a221oi_1
X_4218_ _1049_ _1041_ _1045_ VPWR VGND sg13g2_nand2_1
X_5198_ _1992_ _1991_ _1988_ VPWR VGND sg13g2_nand2b_1
X_4149_ net819 net869 net813 net867 _0984_ VPWR VGND sg13g2_and4_1
XFILLER_44_839 VPWR VGND sg13g2_fill_2
XFILLER_43_305 VPWR VGND sg13g2_fill_2
XFILLER_24_552 VPWR VGND sg13g2_fill_2
Xclkload0 clknet_4_1_0_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_4_968 VPWR VGND sg13g2_decap_8
XFILLER_47_666 VPWR VGND sg13g2_fill_1
XFILLER_42_393 VPWR VGND sg13g2_fill_1
X_3520_ _0381_ _0317_ _0382_ VPWR VGND sg13g2_xor2_1
X_3451_ _0314_ _0306_ _0310_ VPWR VGND sg13g2_nand2_1
X_3382_ net937 net991 net932 net989 _2964_ VPWR VGND sg13g2_and4_1
X_6170_ net1078 VGND VPWR net152 mac1.sum_lvl1_ff\[43\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_5121_ VGND VPWR _1917_ _1915_ _1869_ sg13g2_or2_1
X_5052_ _1847_ _1846_ _1816_ _1850_ VPWR VGND sg13g2_a21o_1
X_4003_ _0845_ _0841_ _0846_ VPWR VGND sg13g2_xor2_1
XFILLER_37_154 VPWR VGND sg13g2_fill_1
XFILLER_38_699 VPWR VGND sg13g2_fill_2
X_5954_ net871 _0228_ VPWR VGND sg13g2_buf_1
X_4905_ _1711_ net872 DP_4.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_5885_ _2567_ VPWR _0225_ VGND net761 _2568_ sg13g2_o21ai_1
XFILLER_21_522 VPWR VGND sg13g2_fill_2
X_4836_ VGND VPWR _1645_ _1643_ _1619_ sg13g2_or2_1
X_4767_ VGND VPWR _1578_ _1576_ _1537_ sg13g2_or2_1
X_3718_ _0539_ _0573_ _0574_ VPWR VGND sg13g2_nor2b_1
X_4698_ _1506_ VPWR _1511_ VGND _1507_ _1509_ sg13g2_o21ai_1
X_6437_ net1093 VGND VPWR net159 mac2.sum_lvl2_ff\[13\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3649_ _0493_ VPWR _0507_ VGND _0483_ _0494_ sg13g2_o21ai_1
XFILLER_1_927 VPWR VGND sg13g2_decap_8
X_6368_ net1094 VGND VPWR _0131_ mac2.products_ff\[81\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_5319_ _2098_ _2101_ _2102_ _2103_ VPWR VGND sg13g2_nor3_1
Xhold23 mac2.sum_lvl1_ff\[51\] VPWR VGND net63 sg13g2_dlygate4sd3_1
X_6299_ net1023 VGND VPWR net501 mac1.sum_lvl3_ff\[8\] clknet_leaf_2_clk sg13g2_dfrbpq_1
Xhold12 mac2.sum_lvl1_ff\[82\] VPWR VGND net52 sg13g2_dlygate4sd3_1
Xhold56 mac1.sum_lvl1_ff\[37\] VPWR VGND net96 sg13g2_dlygate4sd3_1
Xhold34 mac1.sum_lvl2_ff\[46\] VPWR VGND net74 sg13g2_dlygate4sd3_1
Xhold45 mac2.sum_lvl2_ff\[48\] VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold78 mac2.sum_lvl1_ff\[50\] VPWR VGND net118 sg13g2_dlygate4sd3_1
Xhold89 mac1.sum_lvl2_ff\[53\] VPWR VGND net129 sg13g2_dlygate4sd3_1
XFILLER_21_1004 VPWR VGND sg13g2_decap_8
XFILLER_29_644 VPWR VGND sg13g2_fill_2
Xhold67 mac2.sum_lvl1_ff\[11\] VPWR VGND net107 sg13g2_dlygate4sd3_1
XFILLER_17_817 VPWR VGND sg13g2_fill_2
XFILLER_43_124 VPWR VGND sg13g2_decap_4
XFILLER_28_187 VPWR VGND sg13g2_fill_1
XFILLER_43_157 VPWR VGND sg13g2_fill_2
XFILLER_25_850 VPWR VGND sg13g2_decap_8
XFILLER_25_861 VPWR VGND sg13g2_fill_1
XFILLER_40_864 VPWR VGND sg13g2_decap_8
Xfanout1010 net445 net1010 VPWR VGND sg13g2_buf_8
Xfanout1021 net1025 net1021 VPWR VGND sg13g2_buf_8
Xfanout1032 net1034 net1032 VPWR VGND sg13g2_buf_2
Xfanout1043 net1044 net1043 VPWR VGND sg13g2_buf_8
Xfanout1065 net1066 net1065 VPWR VGND sg13g2_buf_8
Xfanout1054 net1056 net1054 VPWR VGND sg13g2_buf_8
Xfanout1098 rst_n net1098 VPWR VGND sg13g2_buf_8
Xfanout1087 net1098 net1087 VPWR VGND sg13g2_buf_8
Xfanout1076 net1077 net1076 VPWR VGND sg13g2_buf_8
XFILLER_48_975 VPWR VGND sg13g2_decap_8
XFILLER_35_647 VPWR VGND sg13g2_fill_1
XFILLER_37_1000 VPWR VGND sg13g2_decap_8
XFILLER_22_308 VPWR VGND sg13g2_fill_1
X_5670_ _2379_ net326 net763 VPWR VGND sg13g2_nand2_1
X_4621_ _1433_ _1434_ _1428_ _1436_ VPWR VGND sg13g2_nand3_1
X_4552_ _0087_ _1355_ _1368_ VPWR VGND sg13g2_xnor2_1
X_4483_ _1307_ _1302_ _1305_ VPWR VGND sg13g2_xnor2_1
X_3503_ _0365_ net978 net939 net982 net933 VPWR VGND sg13g2_a22oi_1
Xhold504 mac2.sum_lvl2_ff\[10\] VPWR VGND net544 sg13g2_dlygate4sd3_1
X_3434_ _0298_ net983 net939 net985 net935 VPWR VGND sg13g2_a22oi_1
X_6222_ net1020 VGND VPWR net164 mac1.sum_lvl2_ff\[49\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_6153_ net1095 VGND VPWR _0258_ DP_4.matrix\[42\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_44_1026 VPWR VGND sg13g2_fill_2
X_3365_ _2937_ _2950_ _2951_ VPWR VGND sg13g2_nor2_1
X_3296_ _2884_ net891 net1006 VPWR VGND sg13g2_nand2_1
X_6084_ net1070 VGND VPWR _0209_ DP_2.matrix\[41\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5104_ _1863_ VPWR _1900_ VGND _1820_ _1864_ sg13g2_o21ai_1
X_5035_ net797 net793 net842 net839 _1833_ VPWR VGND sg13g2_and4_1
XFILLER_39_986 VPWR VGND sg13g2_decap_8
XFILLER_25_102 VPWR VGND sg13g2_fill_1
XFILLER_26_669 VPWR VGND sg13g2_decap_8
X_5937_ net270 _0195_ VPWR VGND sg13g2_buf_1
X_5868_ _2439_ _2441_ _2558_ VPWR VGND sg13g2_and2_1
X_4819_ _1628_ _1607_ _1629_ VPWR VGND sg13g2_nor2b_1
X_5799_ _2502_ _2503_ _2504_ _2505_ VPWR VGND sg13g2_nor3_1
Xoutput24 net24 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_223 VPWR VGND sg13g2_fill_1
XFILLER_45_923 VPWR VGND sg13g2_decap_8
XFILLER_13_853 VPWR VGND sg13g2_fill_2
XFILLER_12_374 VPWR VGND sg13g2_fill_1
XFILLER_40_694 VPWR VGND sg13g2_fill_2
XFILLER_4_551 VPWR VGND sg13g2_fill_1
X_3150_ _2742_ _2698_ _2741_ VPWR VGND sg13g2_xnor2_1
X_3081_ _2675_ net896 net949 VPWR VGND sg13g2_nand2_1
XFILLER_39_249 VPWR VGND sg13g2_fill_2
XFILLER_35_400 VPWR VGND sg13g2_fill_1
XFILLER_36_934 VPWR VGND sg13g2_decap_8
XFILLER_23_628 VPWR VGND sg13g2_decap_4
X_5722_ _2430_ _2417_ _2429_ VPWR VGND sg13g2_nand2b_1
X_3983_ _0826_ _0809_ _0827_ VPWR VGND sg13g2_xor2_1
X_5653_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] _2362_ VPWR VGND sg13g2_nor2_2
X_5584_ _2305_ VPWR _2308_ VGND _2304_ _2306_ sg13g2_o21ai_1
X_4604_ _1419_ _1417_ _1418_ VPWR VGND sg13g2_nand2b_1
Xhold301 mac1.sum_lvl3_ff\[13\] VPWR VGND net341 sg13g2_dlygate4sd3_1
X_4535_ _1353_ _1350_ _1354_ VPWR VGND sg13g2_xor2_1
Xhold312 DP_3.matrix\[44\] VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold334 _2190_ VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold323 DP_3.matrix\[36\] VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold356 DP_3.matrix\[7\] VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold367 _2165_ VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold345 _0025_ VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold378 mac2.sum_lvl3_ff\[5\] VPWR VGND net418 sg13g2_dlygate4sd3_1
X_4466_ VGND VPWR _1241_ _1261_ _1291_ _1263_ sg13g2_a21oi_1
Xfanout803 net804 net803 VPWR VGND sg13g2_buf_8
X_4397_ _1219_ VPWR _1224_ VGND _1221_ _1222_ sg13g2_o21ai_1
X_3417_ _0281_ _0271_ _0282_ VPWR VGND sg13g2_xor2_1
Xhold389 mac1.sum_lvl3_ff\[20\] VPWR VGND net429 sg13g2_dlygate4sd3_1
X_6205_ net1084 VGND VPWR net46 mac1.sum_lvl2_ff\[29\] clknet_leaf_48_clk sg13g2_dfrbpq_2
Xfanout814 net816 net814 VPWR VGND sg13g2_buf_2
Xfanout825 net350 net825 VPWR VGND sg13g2_buf_8
Xfanout858 net860 net858 VPWR VGND sg13g2_buf_8
X_3348_ _2906_ _2932_ _2934_ VPWR VGND sg13g2_and2_1
X_6136_ net1085 VGND VPWR net179 mac1.sum_lvl1_ff\[13\] clknet_leaf_43_clk sg13g2_dfrbpq_1
Xfanout847 DP_3.matrix\[76\] net847 VPWR VGND sg13g2_buf_2
Xfanout836 net837 net836 VPWR VGND sg13g2_buf_1
Xfanout869 net329 net869 VPWR VGND sg13g2_buf_8
X_6067_ net1014 VGND VPWR _0101_ mac1.products_ff\[142\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3279_ _2868_ _2822_ _2866_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_219 VPWR VGND sg13g2_fill_2
XFILLER_26_24 VPWR VGND sg13g2_fill_2
XFILLER_26_411 VPWR VGND sg13g2_fill_2
XFILLER_27_945 VPWR VGND sg13g2_decap_8
X_5018_ _1808_ VPWR _1816_ VGND _1788_ _1809_ sg13g2_o21ai_1
XFILLER_42_959 VPWR VGND sg13g2_decap_8
XFILLER_21_160 VPWR VGND sg13g2_fill_2
XFILLER_42_56 VPWR VGND sg13g2_fill_2
XFILLER_6_838 VPWR VGND sg13g2_decap_8
XFILLER_33_937 VPWR VGND sg13g2_decap_8
XFILLER_34_1003 VPWR VGND sg13g2_decap_8
XFILLER_8_197 VPWR VGND sg13g2_fill_1
X_4320_ _1137_ VPWR _1149_ VGND _1145_ _1147_ sg13g2_o21ai_1
X_4251_ _1073_ VPWR _1081_ VGND _1053_ _1074_ sg13g2_o21ai_1
X_3202_ VGND VPWR _2793_ _2792_ _2745_ sg13g2_or2_1
X_4182_ _1013_ _1012_ _1007_ _1015_ VPWR VGND sg13g2_a21o_1
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
X_3133_ VGND VPWR _2723_ _2724_ _2726_ _2694_ sg13g2_a21oi_1
X_3064_ _2632_ _2656_ _2657_ _2659_ VPWR VGND sg13g2_nor3_1
XFILLER_35_252 VPWR VGND sg13g2_fill_1
XFILLER_35_263 VPWR VGND sg13g2_fill_1
X_3966_ _0779_ VPWR _0810_ VGND _0770_ _0780_ sg13g2_o21ai_1
X_5705_ _2413_ net771 _2412_ net764 net891 VPWR VGND sg13g2_a22oi_1
X_3897_ _0721_ _0740_ _0742_ _0743_ VPWR VGND sg13g2_or3_1
X_5636_ net21 _2346_ _2348_ VPWR VGND sg13g2_xnor2_1
X_5567_ VGND VPWR _2292_ _2294_ _2296_ net399 sg13g2_a21oi_1
X_4518_ VGND VPWR _1323_ _1339_ _1340_ _1338_ sg13g2_a21oi_1
Xhold131 mac1.sum_lvl2_ff\[40\] VPWR VGND net171 sg13g2_dlygate4sd3_1
Xhold153 mac1.sum_lvl1_ff\[79\] VPWR VGND net193 sg13g2_dlygate4sd3_1
Xhold120 mac1.sum_lvl1_ff\[40\] VPWR VGND net160 sg13g2_dlygate4sd3_1
Xhold142 mac2.sum_lvl1_ff\[74\] VPWR VGND net182 sg13g2_dlygate4sd3_1
X_5498_ _2241_ _2242_ _0036_ VPWR VGND sg13g2_nor2b_2
X_4449_ _1254_ VPWR _1274_ VGND _1251_ _1255_ sg13g2_o21ai_1
Xhold164 mac1.products_ff\[4\] VPWR VGND net204 sg13g2_dlygate4sd3_1
Xhold186 mac1.sum_lvl2_ff\[52\] VPWR VGND net226 sg13g2_dlygate4sd3_1
Xhold175 mac1.sum_lvl1_ff\[51\] VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold197 mac1.products_ff\[74\] VPWR VGND net237 sg13g2_dlygate4sd3_1
X_6119_ net1076 VGND VPWR _0232_ DP_3.matrix\[40\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_46_528 VPWR VGND sg13g2_decap_4
XFILLER_46_517 VPWR VGND sg13g2_decap_8
XFILLER_14_425 VPWR VGND sg13g2_fill_1
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_23_970 VPWR VGND sg13g2_decap_8
XFILLER_2_874 VPWR VGND sg13g2_decap_4
XFILLER_49_333 VPWR VGND sg13g2_fill_1
XFILLER_49_366 VPWR VGND sg13g2_fill_2
XFILLER_17_263 VPWR VGND sg13g2_fill_2
X_3820_ _0663_ VPWR _0668_ VGND _0664_ _0666_ sg13g2_o21ai_1
XFILLER_14_992 VPWR VGND sg13g2_decap_8
X_3751_ _0110_ _0588_ _0604_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_462 VPWR VGND sg13g2_fill_1
XFILLER_9_495 VPWR VGND sg13g2_fill_2
X_3682_ VGND VPWR _0539_ _0538_ _0487_ sg13g2_or2_1
X_6470_ net1034 VGND VPWR _0037_ mac2.sum_lvl3_ff\[14\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5421_ net323 mac1.sum_lvl3_ff\[32\] _2183_ VPWR VGND sg13g2_xor2_1
X_5352_ _0003_ _2126_ net536 VPWR VGND sg13g2_xnor2_1
X_4303_ _1132_ net807 net861 VPWR VGND sg13g2_nand2_1
X_5283_ _2072_ _2059_ _2074_ VPWR VGND sg13g2_xor2_1
X_4234_ _1065_ net860 net817 net862 net814 VPWR VGND sg13g2_a22oi_1
X_4165_ _0999_ _0990_ _0997_ VPWR VGND sg13g2_xnor2_1
X_3116_ _2709_ net896 net946 VPWR VGND sg13g2_nand2_1
X_4096_ _0936_ net961 net907 VPWR VGND sg13g2_nand2_1
X_3047_ _2623_ VPWR _2642_ VGND _2621_ _2624_ sg13g2_o21ai_1
X_4998_ _1797_ net791 net847 VPWR VGND sg13g2_nand2_1
X_3949_ _0791_ _0790_ _0792_ _0794_ VPWR VGND sg13g2_a21o_1
XFILLER_20_984 VPWR VGND sg13g2_decap_8
X_5619_ mac1.total_sum\[10\] mac2.total_sum\[10\] _2335_ VPWR VGND sg13g2_and2_1
XFILLER_24_1002 VPWR VGND sg13g2_decap_8
XFILLER_19_506 VPWR VGND sg13g2_fill_1
XFILLER_47_859 VPWR VGND sg13g2_fill_1
XFILLER_46_347 VPWR VGND sg13g2_fill_1
XFILLER_42_597 VPWR VGND sg13g2_fill_2
XFILLER_42_586 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_13_91 VPWR VGND sg13g2_fill_2
XFILLER_7_999 VPWR VGND sg13g2_decap_8
XFILLER_6_465 VPWR VGND sg13g2_fill_1
XFILLER_49_163 VPWR VGND sg13g2_fill_2
XFILLER_37_358 VPWR VGND sg13g2_fill_1
X_5970_ net819 _0252_ VPWR VGND sg13g2_buf_1
X_4921_ _1722_ _1716_ _0091_ VPWR VGND sg13g2_xor2_1
X_4852_ _1659_ _1658_ _1661_ VPWR VGND sg13g2_xor2_1
X_3803_ _0652_ _0650_ _0651_ VPWR VGND sg13g2_nand2_1
X_4783_ _1594_ _1584_ _1593_ VPWR VGND sg13g2_nand2b_1
X_3734_ _0579_ _0581_ _0589_ VPWR VGND sg13g2_and2_1
X_3665_ _0523_ _0518_ _0521_ VPWR VGND sg13g2_xnor2_1
X_6453_ net1097 VGND VPWR net130 mac2.sum_lvl2_ff\[32\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_5404_ mac1.sum_lvl3_ff\[29\] net293 _2169_ VPWR VGND sg13g2_nor2_1
XFILLER_47_1002 VPWR VGND sg13g2_decap_8
X_3596_ _0456_ _0451_ _0455_ VPWR VGND sg13g2_nand2_1
X_6384_ net1032 VGND VPWR _0153_ mac2.products_ff\[149\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5335_ mac1.sum_lvl2_ff\[29\] net548 _2115_ VPWR VGND sg13g2_and2_1
X_5266_ _2030_ _2055_ _2057_ VPWR VGND sg13g2_and2_1
X_4217_ _0127_ _1021_ _1048_ VPWR VGND sg13g2_xnor2_1
X_5197_ _1990_ _1946_ _1991_ VPWR VGND sg13g2_xor2_1
XFILLER_29_837 VPWR VGND sg13g2_fill_1
X_4148_ net871 net811 _0983_ VPWR VGND sg13g2_and2_1
X_4079_ VGND VPWR _0875_ _0880_ _0920_ _0892_ sg13g2_a21oi_1
XFILLER_37_881 VPWR VGND sg13g2_decap_8
XFILLER_11_269 VPWR VGND sg13g2_fill_1
Xclkload1 clknet_4_2_0_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_947 VPWR VGND sg13g2_decap_8
XFILLER_46_144 VPWR VGND sg13g2_fill_2
XFILLER_28_881 VPWR VGND sg13g2_decap_8
XFILLER_34_328 VPWR VGND sg13g2_fill_1
XFILLER_11_770 VPWR VGND sg13g2_fill_1
X_3450_ _0105_ _0286_ _0313_ VPWR VGND sg13g2_xnor2_1
X_3381_ net993 net930 _2963_ VPWR VGND sg13g2_and2_1
X_5120_ _1916_ net789 net841 VPWR VGND sg13g2_nand2_1
XFILLER_3_991 VPWR VGND sg13g2_decap_8
X_5051_ VGND VPWR _1846_ _1847_ _1849_ _1816_ sg13g2_a21oi_1
X_4002_ _0845_ _0802_ _0843_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_829 VPWR VGND sg13g2_fill_1
X_5953_ net888 _0219_ VPWR VGND sg13g2_buf_1
X_4904_ _1698_ VPWR _1710_ VGND _1671_ _1696_ sg13g2_o21ai_1
X_5884_ _2477_ _2458_ _2568_ VPWR VGND sg13g2_xor2_1
XFILLER_34_884 VPWR VGND sg13g2_decap_8
XFILLER_40_309 VPWR VGND sg13g2_fill_1
X_4835_ _1619_ _1643_ _1644_ VPWR VGND sg13g2_nor2_1
X_4766_ _1577_ net879 DP_4.matrix\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_21_589 VPWR VGND sg13g2_fill_1
X_3717_ _0573_ _0568_ _0571_ VPWR VGND sg13g2_xnor2_1
X_4697_ _1506_ _1507_ _1509_ _1510_ VPWR VGND sg13g2_or3_1
X_6436_ net1094 VGND VPWR net238 mac2.sum_lvl2_ff\[12\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3648_ _0480_ _0474_ _0482_ _0506_ VPWR VGND sg13g2_a21o_1
XFILLER_1_906 VPWR VGND sg13g2_decap_8
X_3579_ _0438_ _0434_ _0439_ VPWR VGND sg13g2_xor2_1
X_6367_ net1091 VGND VPWR _0130_ mac2.products_ff\[80\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_5318_ VPWR VGND _2096_ _2095_ _2094_ mac1.sum_lvl2_ff\[24\] _2102_ mac1.sum_lvl2_ff\[5\]
+ sg13g2_a221oi_1
X_6298_ net1023 VGND VPWR _0013_ mac1.sum_lvl3_ff\[7\] clknet_leaf_1_clk sg13g2_dfrbpq_1
Xhold13 mac1.sum_lvl2_ff\[49\] VPWR VGND net53 sg13g2_dlygate4sd3_1
X_5249_ _2040_ _2014_ _2041_ VPWR VGND sg13g2_xor2_1
Xhold24 mac1.products_ff\[5\] VPWR VGND net64 sg13g2_dlygate4sd3_1
Xhold46 mac1.products_ff\[72\] VPWR VGND net86 sg13g2_dlygate4sd3_1
Xhold35 mac1.products_ff\[82\] VPWR VGND net75 sg13g2_dlygate4sd3_1
XFILLER_29_612 VPWR VGND sg13g2_fill_1
Xhold68 mac2.sum_lvl1_ff\[6\] VPWR VGND net108 sg13g2_dlygate4sd3_1
Xhold79 mac2.sum_lvl1_ff\[37\] VPWR VGND net119 sg13g2_dlygate4sd3_1
Xhold57 mac2.products_ff\[148\] VPWR VGND net97 sg13g2_dlygate4sd3_1
XFILLER_25_840 VPWR VGND sg13g2_fill_1
XFILLER_4_777 VPWR VGND sg13g2_fill_2
Xfanout1000 DP_3.matrix\[44\] net1000 VPWR VGND sg13g2_buf_1
Xfanout1022 net1023 net1022 VPWR VGND sg13g2_buf_8
Xfanout1011 DP_1.matrix\[8\] net1011 VPWR VGND sg13g2_buf_1
Xfanout1044 net1045 net1044 VPWR VGND sg13g2_buf_8
XFILLER_0_983 VPWR VGND sg13g2_decap_8
Xfanout1033 net1034 net1033 VPWR VGND sg13g2_buf_8
Xfanout1055 net1056 net1055 VPWR VGND sg13g2_buf_8
XFILLER_48_954 VPWR VGND sg13g2_decap_8
Xfanout1066 net1077 net1066 VPWR VGND sg13g2_buf_8
Xfanout1077 net1098 net1077 VPWR VGND sg13g2_buf_8
Xfanout1088 net1091 net1088 VPWR VGND sg13g2_buf_8
XFILLER_35_637 VPWR VGND sg13g2_fill_2
XFILLER_34_125 VPWR VGND sg13g2_fill_1
XFILLER_34_158 VPWR VGND sg13g2_fill_2
XFILLER_43_692 VPWR VGND sg13g2_fill_1
X_4620_ _1435_ _1428_ _1433_ _1434_ VPWR VGND sg13g2_and3_1
X_4551_ _1355_ _1368_ _1369_ VPWR VGND sg13g2_nor2b_1
X_4482_ _1306_ _1305_ _1302_ VPWR VGND sg13g2_nand2b_1
X_3502_ net933 net981 net938 _0364_ VPWR VGND net978 sg13g2_nand4_1
Xhold505 _2226_ VPWR VGND net545 sg13g2_dlygate4sd3_1
X_3433_ net935 net985 net939 _0297_ VPWR VGND net983 sg13g2_nand4_1
X_6221_ net1019 VGND VPWR net207 mac1.sum_lvl2_ff\[48\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_6152_ net1092 VGND VPWR _0257_ DP_4.matrix\[41\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_44_1005 VPWR VGND sg13g2_decap_8
X_3364_ _2948_ _2938_ _2950_ VPWR VGND sg13g2_xor2_1
X_5103_ _0158_ _1854_ _1898_ VPWR VGND sg13g2_xnor2_1
X_3295_ _2883_ net1007 net893 net943 net890 VPWR VGND sg13g2_a22oi_1
X_6083_ net1081 VGND VPWR _0208_ DP_2.matrix\[40\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_5034_ _1832_ net791 net845 VPWR VGND sg13g2_nand2_1
XFILLER_38_442 VPWR VGND sg13g2_fill_2
XFILLER_39_965 VPWR VGND sg13g2_decap_8
X_5936_ net278 _0194_ VPWR VGND sg13g2_buf_1
X_5867_ _2557_ net925 net755 VPWR VGND sg13g2_nand2b_1
XFILLER_22_876 VPWR VGND sg13g2_fill_2
X_4818_ _1628_ _1608_ _1627_ VPWR VGND sg13g2_xnor2_1
X_5798_ net796 net767 _2504_ VPWR VGND sg13g2_nor2_1
X_4749_ _1560_ _1543_ _1561_ VPWR VGND sg13g2_xor2_1
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
X_6419_ net1027 VGND VPWR net1 DP_1.I_range.out_data\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_2
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_45_902 VPWR VGND sg13g2_decap_8
XFILLER_45_979 VPWR VGND sg13g2_decap_8
XFILLER_16_147 VPWR VGND sg13g2_fill_2
X_3080_ _2645_ VPWR _2674_ VGND _2643_ _2646_ sg13g2_o21ai_1
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_36_913 VPWR VGND sg13g2_decap_8
X_3982_ _0826_ _0810_ _0824_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_489 VPWR VGND sg13g2_fill_2
X_5721_ _2428_ _2425_ _2424_ _2429_ VPWR VGND sg13g2_a21o_1
XFILLER_15_180 VPWR VGND sg13g2_fill_2
X_5652_ _2361_ DP_1.Q_range.out_data\[5\] DP_1.Q_range.out_data\[6\] VPWR VGND sg13g2_nand2b_1
XFILLER_30_172 VPWR VGND sg13g2_decap_4
XFILLER_31_695 VPWR VGND sg13g2_fill_2
X_5583_ net26 _2304_ _2307_ VPWR VGND sg13g2_xnor2_1
X_4603_ _1418_ DP_3.matrix\[0\] net821 VPWR VGND sg13g2_nand2_1
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
Xhold302 _2187_ VPWR VGND net342 sg13g2_dlygate4sd3_1
X_4534_ _1351_ _1352_ _1353_ VPWR VGND sg13g2_nor2_1
Xhold324 DP_3.matrix\[5\] VPWR VGND net364 sg13g2_dlygate4sd3_1
XFILLER_7_390 VPWR VGND sg13g2_fill_1
Xhold313 mac1.sum_lvl3_ff\[4\] VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold335 _0021_ VPWR VGND net375 sg13g2_dlygate4sd3_1
Xhold357 _2571_ VPWR VGND net397 sg13g2_dlygate4sd3_1
Xhold346 DP_3.matrix\[6\] VPWR VGND net386 sg13g2_dlygate4sd3_1
X_4465_ _1290_ _1269_ _1289_ VPWR VGND sg13g2_xnor2_1
Xhold368 _0030_ VPWR VGND net408 sg13g2_dlygate4sd3_1
Xfanout804 net467 net804 VPWR VGND sg13g2_buf_8
X_4396_ _1219_ _1221_ _1222_ _1223_ VPWR VGND sg13g2_nor3_1
X_3416_ _0281_ _0279_ _0280_ VPWR VGND sg13g2_nand2_1
X_6204_ net1081 VGND VPWR net239 mac1.sum_lvl2_ff\[28\] clknet_leaf_49_clk sg13g2_dfrbpq_2
Xhold379 _2264_ VPWR VGND net419 sg13g2_dlygate4sd3_1
Xfanout815 net816 net815 VPWR VGND sg13g2_buf_1
X_6135_ net1061 VGND VPWR _0243_ DP_3.matrix\[79\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3347_ _2933_ _2932_ _0098_ VPWR VGND sg13g2_xor2_1
Xfanout837 net376 net837 VPWR VGND sg13g2_buf_1
Xfanout848 DP_3.matrix\[75\] net848 VPWR VGND sg13g2_buf_8
Xfanout826 DP_4.matrix\[3\] net826 VPWR VGND sg13g2_buf_1
Xfanout859 net860 net859 VPWR VGND sg13g2_buf_1
X_6066_ net1044 VGND VPWR _0197_ DP_2.matrix\[1\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3278_ VGND VPWR _2867_ _2865_ _2823_ sg13g2_or2_1
X_5017_ _1815_ _1814_ _0156_ VPWR VGND sg13g2_xor2_1
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_39_773 VPWR VGND sg13g2_decap_8
XFILLER_42_938 VPWR VGND sg13g2_decap_8
XFILLER_13_139 VPWR VGND sg13g2_fill_1
X_5919_ net997 _0168_ VPWR VGND sg13g2_buf_1
XFILLER_22_640 VPWR VGND sg13g2_fill_2
XFILLER_22_651 VPWR VGND sg13g2_decap_8
XFILLER_10_857 VPWR VGND sg13g2_fill_2
XFILLER_10_846 VPWR VGND sg13g2_fill_2
XFILLER_5_338 VPWR VGND sg13g2_fill_1
XFILLER_49_515 VPWR VGND sg13g2_decap_4
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_559 VPWR VGND sg13g2_fill_1
XFILLER_36_209 VPWR VGND sg13g2_fill_1
XFILLER_33_916 VPWR VGND sg13g2_decap_8
XFILLER_12_150 VPWR VGND sg13g2_decap_8
XFILLER_12_161 VPWR VGND sg13g2_fill_1
XFILLER_12_172 VPWR VGND sg13g2_fill_2
XFILLER_8_154 VPWR VGND sg13g2_fill_2
XFILLER_8_187 VPWR VGND sg13g2_fill_2
XFILLER_4_382 VPWR VGND sg13g2_fill_2
X_4250_ _1080_ _1079_ _0134_ VPWR VGND sg13g2_xor2_1
X_3201_ _2792_ net894 net944 VPWR VGND sg13g2_nand2_1
X_4181_ _1012_ _1013_ _1007_ _1014_ VPWR VGND sg13g2_nand3_1
X_3132_ _2723_ _2724_ _2694_ _2725_ VPWR VGND sg13g2_nand3_1
X_3063_ _2654_ _2655_ _2618_ _2658_ VPWR VGND sg13g2_nand3_1
XFILLER_36_710 VPWR VGND sg13g2_fill_1
XFILLER_48_592 VPWR VGND sg13g2_decap_8
XFILLER_24_916 VPWR VGND sg13g2_fill_2
X_3965_ _0807_ _0799_ _0809_ VPWR VGND sg13g2_xor2_1
X_3896_ VGND VPWR _0738_ _0739_ _0742_ _0722_ sg13g2_a21oi_1
X_5704_ net927 net911 net775 _2412_ VPWR VGND sg13g2_mux2_1
X_5635_ _2348_ VPWR _2349_ VGND _2344_ _2345_ sg13g2_o21ai_1
Xhold110 mac1.products_ff\[12\] VPWR VGND net150 sg13g2_dlygate4sd3_1
X_5566_ _2295_ mac2.sum_lvl3_ff\[33\] net398 VPWR VGND sg13g2_xnor2_1
X_4517_ _1339_ _1323_ _0132_ VPWR VGND sg13g2_xor2_1
Xhold143 mac1.sum_lvl1_ff\[42\] VPWR VGND net183 sg13g2_dlygate4sd3_1
Xhold132 mac1.sum_lvl1_ff\[76\] VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold121 mac1.products_ff\[139\] VPWR VGND net161 sg13g2_dlygate4sd3_1
X_5497_ _2239_ _2240_ net512 _2242_ VPWR VGND sg13g2_nand3_1
X_4448_ _1273_ _1272_ _1270_ VPWR VGND sg13g2_nand2b_1
Xhold165 mac1.sum_lvl1_ff\[1\] VPWR VGND net205 sg13g2_dlygate4sd3_1
Xhold176 mac1.sum_lvl1_ff\[80\] VPWR VGND net216 sg13g2_dlygate4sd3_1
Xhold154 mac2.sum_lvl1_ff\[77\] VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold198 mac2.sum_lvl1_ff\[12\] VPWR VGND net238 sg13g2_dlygate4sd3_1
Xhold187 mac2.sum_lvl1_ff\[8\] VPWR VGND net227 sg13g2_dlygate4sd3_1
X_4379_ _1171_ VPWR _1206_ VGND _1168_ _1172_ sg13g2_o21ai_1
X_6118_ net1068 VGND VPWR net230 mac1.sum_lvl1_ff\[7\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_6049_ net1039 VGND VPWR _0064_ mac1.products_ff\[136\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_2_1013 VPWR VGND sg13g2_decap_8
XFILLER_15_938 VPWR VGND sg13g2_decap_8
XFILLER_41_212 VPWR VGND sg13g2_fill_2
XFILLER_5_179 VPWR VGND sg13g2_fill_1
XFILLER_33_702 VPWR VGND sg13g2_fill_1
XFILLER_33_713 VPWR VGND sg13g2_fill_2
XFILLER_13_470 VPWR VGND sg13g2_fill_1
XFILLER_14_971 VPWR VGND sg13g2_decap_8
X_3750_ VPWR _0605_ _0604_ VGND sg13g2_inv_1
X_3681_ _0538_ DP_2.matrix\[5\] net1011 VPWR VGND sg13g2_nand2_1
X_5420_ mac1.sum_lvl3_ff\[32\] net323 _2182_ VPWR VGND sg13g2_nor2_1
X_5351_ _2128_ VPWR _2129_ VGND _2124_ _2125_ sg13g2_o21ai_1
X_5282_ VGND VPWR _2073_ _2072_ _2059_ sg13g2_or2_1
X_4302_ _1131_ net866 net805 VPWR VGND sg13g2_nand2_1
XFILLER_4_190 VPWR VGND sg13g2_fill_2
X_4233_ net814 net862 net817 _1064_ VPWR VGND net860 sg13g2_nand4_1
X_4164_ _0998_ _0997_ _0990_ VPWR VGND sg13g2_nand2b_1
X_3115_ _2677_ VPWR _2708_ VGND _2675_ _2678_ sg13g2_o21ai_1
X_4095_ _0935_ net966 net1004 VPWR VGND sg13g2_nand2_1
X_3046_ _2639_ _2636_ _2641_ VPWR VGND sg13g2_xor2_1
XFILLER_36_551 VPWR VGND sg13g2_fill_1
XFILLER_12_919 VPWR VGND sg13g2_fill_1
XFILLER_11_418 VPWR VGND sg13g2_fill_1
XFILLER_17_1010 VPWR VGND sg13g2_decap_8
X_4997_ _1767_ VPWR _1796_ VGND _1765_ _1768_ sg13g2_o21ai_1
X_3948_ _0791_ _0792_ _0790_ _0793_ VPWR VGND sg13g2_nand3_1
X_3879_ VGND VPWR _0725_ _0724_ _0689_ sg13g2_or2_1
X_5618_ net18 _2332_ _2334_ VPWR VGND sg13g2_xnor2_1
X_5549_ mac2.sum_lvl3_ff\[10\] net380 _2281_ VPWR VGND sg13g2_xor2_1
XFILLER_2_105 VPWR VGND sg13g2_fill_2
XFILLER_48_78 VPWR VGND sg13g2_fill_2
XFILLER_46_326 VPWR VGND sg13g2_fill_2
XFILLER_27_540 VPWR VGND sg13g2_fill_1
XFILLER_30_749 VPWR VGND sg13g2_decap_8
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_31_1018 VPWR VGND sg13g2_decap_8
XFILLER_10_484 VPWR VGND sg13g2_decap_8
XFILLER_7_978 VPWR VGND sg13g2_decap_8
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_37_304 VPWR VGND sg13g2_fill_2
XFILLER_18_562 VPWR VGND sg13g2_decap_8
XFILLER_46_882 VPWR VGND sg13g2_decap_8
X_4920_ _1723_ _1716_ _1722_ VPWR VGND sg13g2_nand2_1
X_4851_ VGND VPWR _1660_ _1659_ _1658_ sg13g2_or2_1
X_3802_ _0651_ _0631_ _0633_ VPWR VGND sg13g2_nand2_1
X_4782_ _1593_ _1585_ _1592_ VPWR VGND sg13g2_xnor2_1
X_3733_ VPWR VGND _0564_ _0584_ _0587_ _0559_ _0588_ _0583_ sg13g2_a221oi_1
X_3664_ _0522_ _0521_ _0518_ VPWR VGND sg13g2_nand2b_1
X_6452_ net1096 VGND VPWR net141 mac2.sum_lvl2_ff\[31\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_5403_ _2168_ mac1.sum_lvl3_ff\[29\] net293 VPWR VGND sg13g2_nand2_1
X_3595_ _0453_ _0454_ _0455_ VPWR VGND sg13g2_nor2_1
X_6383_ net1033 VGND VPWR _0152_ mac2.products_ff\[148\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_5334_ _0015_ _2112_ net547 VPWR VGND sg13g2_xnor2_1
X_5265_ _0153_ _2055_ _2056_ VPWR VGND sg13g2_xnor2_1
X_5196_ _1990_ net844 net784 VPWR VGND sg13g2_nand2_1
X_4216_ _1048_ _1047_ _1046_ VPWR VGND sg13g2_nand2b_1
X_4147_ _0981_ _0982_ _0080_ VPWR VGND sg13g2_nor2_1
X_4078_ _0917_ _0905_ _0919_ VPWR VGND sg13g2_xor2_1
XFILLER_37_860 VPWR VGND sg13g2_decap_8
X_3029_ _2621_ _2622_ _2624_ _2625_ VPWR VGND sg13g2_or3_1
Xclkload2 clknet_4_3_0_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_4_926 VPWR VGND sg13g2_decap_8
XFILLER_28_860 VPWR VGND sg13g2_decap_8
XFILLER_43_885 VPWR VGND sg13g2_decap_8
X_3380_ _2961_ _2962_ _0070_ VPWR VGND sg13g2_nor2_1
XFILLER_3_970 VPWR VGND sg13g2_decap_8
X_5050_ _1846_ _1847_ _1816_ _1848_ VPWR VGND sg13g2_nand3_1
X_4001_ VGND VPWR _0844_ _0842_ _0803_ sg13g2_or2_1
X_5952_ net280 _0218_ VPWR VGND sg13g2_buf_1
XFILLER_37_167 VPWR VGND sg13g2_decap_4
X_4903_ VGND VPWR _1679_ _1702_ _1709_ _1704_ sg13g2_a21oi_1
X_5883_ _2567_ net876 net761 VPWR VGND sg13g2_nand2_1
XFILLER_21_513 VPWR VGND sg13g2_fill_1
X_4834_ _1643_ net875 DP_4.matrix\[7\] VPWR VGND sg13g2_nand2_2
XFILLER_21_524 VPWR VGND sg13g2_fill_1
X_4765_ _1576_ net879 net820 VPWR VGND sg13g2_nand2_1
XFILLER_14_1013 VPWR VGND sg13g2_decap_8
X_3716_ _0572_ _0571_ _0568_ VPWR VGND sg13g2_nand2b_1
X_4696_ _1509_ net1001 net835 net873 net831 VPWR VGND sg13g2_a22oi_1
X_3647_ _0505_ _0502_ _0106_ VPWR VGND sg13g2_xor2_1
X_6435_ net1096 VGND VPWR net107 mac2.sum_lvl2_ff\[11\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3578_ _0438_ _0388_ _0436_ VPWR VGND sg13g2_xnor2_1
X_6366_ net1088 VGND VPWR _0129_ mac2.products_ff\[79\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_5317_ _2101_ mac1.sum_lvl2_ff\[25\] net514 VPWR VGND sg13g2_xnor2_1
X_6297_ net1023 VGND VPWR _0012_ mac1.sum_lvl3_ff\[6\] clknet_leaf_0_clk sg13g2_dfrbpq_1
Xhold14 mac2.products_ff\[145\] VPWR VGND net54 sg13g2_dlygate4sd3_1
X_5248_ _2040_ net783 net838 VPWR VGND sg13g2_nand2_1
Xhold47 mac1.sum_lvl1_ff\[75\] VPWR VGND net87 sg13g2_dlygate4sd3_1
Xhold25 mac1.products_ff\[9\] VPWR VGND net65 sg13g2_dlygate4sd3_1
Xhold36 mac1.products_ff\[14\] VPWR VGND net76 sg13g2_dlygate4sd3_1
Xhold58 mac1.products_ff\[10\] VPWR VGND net98 sg13g2_dlygate4sd3_1
Xhold69 mac2.sum_lvl1_ff\[3\] VPWR VGND net109 sg13g2_dlygate4sd3_1
X_5179_ VGND VPWR _1896_ _1937_ _1974_ _1938_ sg13g2_a21oi_1
XFILLER_43_159 VPWR VGND sg13g2_fill_1
XFILLER_25_830 VPWR VGND sg13g2_fill_1
XFILLER_25_896 VPWR VGND sg13g2_decap_8
XFILLER_40_899 VPWR VGND sg13g2_decap_8
XFILLER_3_200 VPWR VGND sg13g2_fill_2
XFILLER_4_789 VPWR VGND sg13g2_fill_2
Xfanout1001 net441 net1001 VPWR VGND sg13g2_buf_8
Xfanout1012 net1013 net1012 VPWR VGND sg13g2_buf_8
Xfanout1045 net1048 net1045 VPWR VGND sg13g2_buf_8
Xfanout1023 net1024 net1023 VPWR VGND sg13g2_buf_8
XFILLER_0_962 VPWR VGND sg13g2_decap_8
Xfanout1056 net1063 net1056 VPWR VGND sg13g2_buf_8
Xfanout1034 net1038 net1034 VPWR VGND sg13g2_buf_8
XFILLER_48_933 VPWR VGND sg13g2_decap_8
Xfanout1067 net1069 net1067 VPWR VGND sg13g2_buf_8
Xfanout1078 net1079 net1078 VPWR VGND sg13g2_buf_8
Xfanout1089 net1090 net1089 VPWR VGND sg13g2_buf_8
XFILLER_47_443 VPWR VGND sg13g2_fill_2
XFILLER_19_134 VPWR VGND sg13g2_fill_1
XFILLER_35_605 VPWR VGND sg13g2_fill_2
XFILLER_31_899 VPWR VGND sg13g2_decap_8
X_4550_ _1368_ _1356_ _1366_ VPWR VGND sg13g2_xnor2_1
X_4481_ _1304_ _1277_ _1305_ VPWR VGND sg13g2_xor2_1
X_3501_ net938 net933 net981 net978 _0363_ VPWR VGND sg13g2_and4_1
Xhold506 mac1.sum_lvl2_ff\[9\] VPWR VGND net546 sg13g2_dlygate4sd3_1
X_3432_ net939 net935 net985 net983 _0296_ VPWR VGND sg13g2_and4_1
X_6220_ net1019 VGND VPWR net180 mac1.sum_lvl2_ff\[47\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3363_ _2948_ _2938_ _2949_ VPWR VGND sg13g2_nor2b_1
X_6151_ net1074 VGND VPWR _0256_ DP_4.matrix\[40\] clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
X_5102_ _1853_ _1898_ _1852_ _1899_ VPWR VGND sg13g2_nand3_1
X_3294_ _2869_ _2863_ _2871_ _2882_ VPWR VGND sg13g2_a21o_1
X_6082_ net1019 VGND VPWR _0096_ mac1.products_ff\[147\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_39_944 VPWR VGND sg13g2_decap_8
X_5033_ _1799_ VPWR _1831_ VGND _1797_ _1800_ sg13g2_o21ai_1
X_5935_ net948 _0193_ VPWR VGND sg13g2_buf_1
XFILLER_15_27 VPWR VGND sg13g2_fill_2
XFILLER_25_159 VPWR VGND sg13g2_fill_2
X_5866_ VGND VPWR net755 _2556_ _0202_ _2555_ sg13g2_a21oi_1
X_4817_ _1625_ _1615_ _1627_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_60_clk clknet_4_2_0_clk clknet_leaf_60_clk VPWR VGND sg13g2_buf_8
X_5797_ VGND VPWR net813 net767 _2503_ net780 sg13g2_a21oi_1
X_4748_ _1560_ _1544_ _1558_ VPWR VGND sg13g2_xnor2_1
X_4679_ _1492_ _1491_ _1488_ VPWR VGND sg13g2_nand2b_1
X_6418_ net1094 VGND VPWR net168 mac2.sum_lvl1_ff\[51\] clknet_leaf_35_clk sg13g2_dfrbpq_1
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_737 VPWR VGND sg13g2_fill_1
X_6349_ net1090 VGND VPWR _0139_ mac2.products_ff\[10\] clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_44_413 VPWR VGND sg13g2_fill_1
XFILLER_29_498 VPWR VGND sg13g2_fill_1
XFILLER_45_958 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_51_clk clknet_4_10_0_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
XFILLER_13_855 VPWR VGND sg13g2_fill_1
XFILLER_40_696 VPWR VGND sg13g2_fill_1
XFILLER_8_369 VPWR VGND sg13g2_fill_2
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_39_218 VPWR VGND sg13g2_fill_2
XFILLER_36_969 VPWR VGND sg13g2_decap_8
X_3981_ _0825_ _0810_ _0824_ VPWR VGND sg13g2_nand2_1
XFILLER_23_608 VPWR VGND sg13g2_fill_2
XFILLER_44_991 VPWR VGND sg13g2_decap_8
X_5720_ _2427_ VPWR _2428_ VGND net930 net776 sg13g2_o21ai_1
XFILLER_22_129 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_42_clk clknet_4_12_0_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
X_5651_ _2360_ DP_1.I_range.out_data\[5\] _2359_ VPWR VGND sg13g2_nand2_1
X_5582_ mac2.total_sum\[1\] mac1.total_sum\[1\] _2307_ VPWR VGND sg13g2_xor2_1
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
X_4602_ _1394_ VPWR _1417_ VGND _1371_ _1392_ sg13g2_o21ai_1
X_4533_ _1352_ net882 net833 net829 net884 VPWR VGND sg13g2_a22oi_1
Xhold314 _2151_ VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold303 _0020_ VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold325 DP_3.matrix\[0\] VPWR VGND net365 sg13g2_dlygate4sd3_1
X_4464_ _1289_ _1286_ _1287_ VPWR VGND sg13g2_xnor2_1
X_6203_ net1080 VGND VPWR net192 mac1.sum_lvl2_ff\[27\] clknet_leaf_44_clk sg13g2_dfrbpq_1
Xhold347 DP_2.matrix\[7\] VPWR VGND net387 sg13g2_dlygate4sd3_1
Xhold369 mac1.sum_lvl3_ff\[35\] VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold358 mac2.sum_lvl3_ff\[13\] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold336 DP_4.matrix\[0\] VPWR VGND net376 sg13g2_dlygate4sd3_1
X_4395_ _1222_ net856 net810 net859 net807 VPWR VGND sg13g2_a22oi_1
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_8
X_3415_ _0278_ _0277_ _0272_ _0280_ VPWR VGND sg13g2_a21o_1
Xfanout816 DP_4.matrix\[37\] net816 VPWR VGND sg13g2_buf_2
Xfanout838 net840 net838 VPWR VGND sg13g2_buf_8
X_6134_ net1054 VGND VPWR _0242_ DP_3.matrix\[78\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3346_ _2933_ _2905_ _2911_ VPWR VGND sg13g2_nand2_1
Xfanout827 net366 net827 VPWR VGND sg13g2_buf_8
Xfanout849 net421 net849 VPWR VGND sg13g2_buf_1
X_6065_ net1044 VGND VPWR _0196_ DP_2.matrix\[0\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3277_ _2866_ net947 net889 VPWR VGND sg13g2_nand2_1
XFILLER_27_903 VPWR VGND sg13g2_decap_8
X_5016_ VGND VPWR _1756_ _1782_ _1815_ _1781_ sg13g2_a21oi_1
XFILLER_42_917 VPWR VGND sg13g2_decap_8
X_5918_ net999 _0167_ VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_33_clk clknet_4_13_0_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_5849_ _2423_ _2419_ _2545_ VPWR VGND sg13g2_xor2_1
XFILLER_21_162 VPWR VGND sg13g2_fill_1
XFILLER_42_47 VPWR VGND sg13g2_fill_1
XFILLER_42_58 VPWR VGND sg13g2_fill_1
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_424 VPWR VGND sg13g2_fill_2
XFILLER_18_969 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_4_7_0_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_41_983 VPWR VGND sg13g2_decap_8
XFILLER_8_177 VPWR VGND sg13g2_fill_1
X_3200_ _2791_ net950 net890 VPWR VGND sg13g2_nand2_1
X_4180_ _1008_ VPWR _1013_ VGND _1009_ _1011_ sg13g2_o21ai_1
X_3131_ _2701_ VPWR _2724_ VGND _2720_ _2722_ sg13g2_o21ai_1
X_3062_ _2657_ _2618_ _2654_ _2655_ VPWR VGND sg13g2_and3_1
XFILLER_35_232 VPWR VGND sg13g2_fill_2
X_3964_ _0807_ _0799_ _0808_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_15_clk clknet_4_4_0_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_3895_ _0738_ _0739_ _0722_ _0741_ VPWR VGND sg13g2_nand3_1
X_5703_ net764 net275 _2410_ _2411_ VPWR VGND sg13g2_a21o_1
XFILLER_32_983 VPWR VGND sg13g2_decap_8
X_5634_ mac2.total_sum\[12\] mac1.total_sum\[12\] _2348_ VPWR VGND sg13g2_xor2_1
X_5565_ _0051_ _2291_ net312 VPWR VGND sg13g2_xnor2_1
Xhold100 mac2.sum_lvl1_ff\[5\] VPWR VGND net140 sg13g2_dlygate4sd3_1
X_4516_ _1337_ _1324_ _1339_ VPWR VGND sg13g2_xor2_1
Xhold122 mac1.sum_lvl1_ff\[6\] VPWR VGND net162 sg13g2_dlygate4sd3_1
Xhold133 mac1.sum_lvl1_ff\[43\] VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold111 mac1.sum_lvl1_ff\[8\] VPWR VGND net151 sg13g2_dlygate4sd3_1
Xhold144 mac2.products_ff\[10\] VPWR VGND net184 sg13g2_dlygate4sd3_1
X_5496_ VGND VPWR net512 _2239_ _2241_ _2240_ sg13g2_a21oi_1
X_4447_ VGND VPWR _1272_ _1271_ _1220_ sg13g2_or2_1
Xhold166 mac1.products_ff\[150\] VPWR VGND net206 sg13g2_dlygate4sd3_1
Xhold177 mac1.sum_lvl1_ff\[50\] VPWR VGND net217 sg13g2_dlygate4sd3_1
Xhold155 mac2.products_ff\[4\] VPWR VGND net195 sg13g2_dlygate4sd3_1
Xhold199 mac1.sum_lvl1_ff\[45\] VPWR VGND net239 sg13g2_dlygate4sd3_1
Xhold188 mac2.products_ff\[9\] VPWR VGND net228 sg13g2_dlygate4sd3_1
X_4378_ _1192_ VPWR _1205_ VGND _1176_ _1193_ sg13g2_o21ai_1
X_6117_ net1074 VGND VPWR _0231_ DP_3.matrix\[39\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3329_ _2916_ net943 net887 VPWR VGND sg13g2_nand2_1
X_6048_ net1086 VGND VPWR _0185_ DP_1.matrix\[41\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_41_257 VPWR VGND sg13g2_fill_1
XFILLER_2_821 VPWR VGND sg13g2_fill_2
XFILLER_33_747 VPWR VGND sg13g2_fill_1
XFILLER_14_950 VPWR VGND sg13g2_decap_8
X_3680_ _0537_ net1011 DP_2.matrix\[4\] net980 DP_2.matrix\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_9_497 VPWR VGND sg13g2_fill_1
X_5350_ net535 mac1.sum_lvl2_ff\[31\] _2128_ VPWR VGND sg13g2_xor2_1
X_5281_ _2070_ _2060_ _2072_ VPWR VGND sg13g2_xor2_1
X_4301_ _1103_ VPWR _1130_ VGND _1094_ _1104_ sg13g2_o21ai_1
X_4232_ net817 net814 net862 net860 _1063_ VPWR VGND sg13g2_and4_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ _0995_ _0996_ _0997_ VPWR VGND sg13g2_nor2b_1
X_3114_ _2707_ _2703_ _2706_ VPWR VGND sg13g2_xnor2_1
X_4094_ _0911_ VPWR _0934_ VGND _0908_ _0912_ sg13g2_o21ai_1
XFILLER_49_891 VPWR VGND sg13g2_decap_8
X_3045_ _2640_ _2639_ _2636_ VPWR VGND sg13g2_nand2b_1
X_4996_ _1795_ _1790_ _1793_ VPWR VGND sg13g2_xnor2_1
X_3947_ _0745_ VPWR _0792_ VGND _0685_ _0746_ sg13g2_o21ai_1
X_3878_ _0724_ net914 net968 VPWR VGND sg13g2_nand2_1
X_5617_ mac2.total_sum\[9\] mac1.total_sum\[9\] _2334_ VPWR VGND sg13g2_xor2_1
X_5548_ net380 mac2.sum_lvl3_ff\[10\] _2280_ VPWR VGND sg13g2_and2_1
XFILLER_3_629 VPWR VGND sg13g2_fill_1
X_5479_ VPWR VGND mac2.sum_lvl2_ff\[9\] _2220_ mac2.sum_lvl2_ff\[28\] mac2.sum_lvl2_ff\[27\]
+ _2227_ mac2.sum_lvl2_ff\[8\] sg13g2_a221oi_1
XFILLER_47_817 VPWR VGND sg13g2_decap_8
XFILLER_46_316 VPWR VGND sg13g2_fill_1
XFILLER_11_942 VPWR VGND sg13g2_decap_8
XFILLER_7_957 VPWR VGND sg13g2_decap_8
XFILLER_6_434 VPWR VGND sg13g2_fill_2
XFILLER_1_183 VPWR VGND sg13g2_fill_2
XFILLER_49_165 VPWR VGND sg13g2_fill_1
XFILLER_46_850 VPWR VGND sg13g2_fill_1
XFILLER_33_511 VPWR VGND sg13g2_fill_2
X_4850_ VGND VPWR _1608_ _1627_ _1659_ _1629_ sg13g2_a21oi_1
X_3801_ _0649_ _0639_ _0650_ VPWR VGND sg13g2_xor2_1
X_4781_ _1590_ _1591_ _1592_ VPWR VGND sg13g2_nor2b_1
X_3732_ _0560_ _0585_ _0587_ VPWR VGND sg13g2_and2_1
Xclkload20 clkload20/Y clknet_leaf_49_clk VPWR VGND sg13g2_inv_2
X_3663_ _0520_ _0476_ _0521_ VPWR VGND sg13g2_xor2_1
X_6451_ net1089 VGND VPWR net59 mac2.sum_lvl2_ff\[30\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_5402_ VGND VPWR mac1.sum_lvl3_ff\[28\] mac1.sum_lvl3_ff\[8\] _2167_ _2165_ sg13g2_a21oi_1
X_6382_ net1026 VGND VPWR _0151_ mac2.products_ff\[147\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5333_ net546 mac1.sum_lvl2_ff\[28\] _2114_ VPWR VGND sg13g2_xor2_1
X_3594_ _0454_ net1010 net934 net978 net930 VPWR VGND sg13g2_a22oi_1
X_5264_ VGND VPWR _2030_ _2034_ _2056_ _2029_ sg13g2_a21oi_1
X_5195_ _1989_ net844 net781 VPWR VGND sg13g2_nand2_1
X_4215_ _1019_ VPWR _1047_ VGND _1043_ _1044_ sg13g2_o21ai_1
X_4146_ _0982_ net813 net871 net869 net819 VPWR VGND sg13g2_a22oi_1
X_4077_ VGND VPWR _0918_ _0917_ _0905_ sg13g2_or2_1
X_3028_ _2624_ net949 net904 net952 net898 VPWR VGND sg13g2_a22oi_1
XFILLER_24_522 VPWR VGND sg13g2_decap_8
XFILLER_24_588 VPWR VGND sg13g2_fill_2
X_4979_ _1779_ _1740_ _1776_ _1777_ VPWR VGND sg13g2_and3_1
XFILLER_11_249 VPWR VGND sg13g2_fill_1
XFILLER_20_750 VPWR VGND sg13g2_fill_1
Xclkload3 clknet_4_5_0_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_47_603 VPWR VGND sg13g2_decap_8
XFILLER_46_146 VPWR VGND sg13g2_fill_1
XFILLER_30_503 VPWR VGND sg13g2_fill_1
XFILLER_30_569 VPWR VGND sg13g2_decap_4
X_4000_ _0843_ net968 net908 VPWR VGND sg13g2_nand2_1
XFILLER_1_41 VPWR VGND sg13g2_fill_1
X_5951_ net891 _0217_ VPWR VGND sg13g2_buf_1
XFILLER_25_319 VPWR VGND sg13g2_fill_2
X_4902_ VGND VPWR _1691_ _1707_ _1708_ _1706_ sg13g2_a21oi_1
X_5882_ _2565_ VPWR _0224_ VGND net759 _2566_ sg13g2_o21ai_1
X_4833_ _1642_ DP_3.matrix\[4\] net996 VPWR VGND sg13g2_nand2_1
XFILLER_33_385 VPWR VGND sg13g2_fill_2
X_4764_ _1575_ net883 net996 VPWR VGND sg13g2_nand2_1
X_3715_ _0570_ _0544_ _0571_ VPWR VGND sg13g2_xor2_1
X_6434_ net1096 VGND VPWR net50 mac2.sum_lvl2_ff\[10\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_4695_ net831 net873 net836 _1508_ VPWR VGND net1001 sg13g2_nand4_1
X_3646_ _0505_ _0503_ _0504_ VPWR VGND sg13g2_nand2b_1
X_3577_ VGND VPWR _0437_ _0435_ _0389_ sg13g2_or2_1
X_6365_ net1088 VGND VPWR _0128_ mac2.products_ff\[78\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5316_ mac1.sum_lvl2_ff\[25\] mac1.sum_lvl2_ff\[6\] _2100_ VPWR VGND sg13g2_and2_1
X_6296_ net1023 VGND VPWR _0011_ mac1.sum_lvl3_ff\[5\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5247_ _2039_ net838 net781 VPWR VGND sg13g2_nand2_1
Xhold15 mac1.sum_lvl2_ff\[50\] VPWR VGND net55 sg13g2_dlygate4sd3_1
Xhold26 mac2.products_ff\[137\] VPWR VGND net66 sg13g2_dlygate4sd3_1
Xhold37 mac2.products_ff\[136\] VPWR VGND net77 sg13g2_dlygate4sd3_1
Xhold59 mac1.products_ff\[11\] VPWR VGND net99 sg13g2_dlygate4sd3_1
XFILLER_21_1018 VPWR VGND sg13g2_decap_8
Xhold48 mac2.sum_lvl1_ff\[44\] VPWR VGND net88 sg13g2_dlygate4sd3_1
X_5178_ _1853_ _1898_ _1852_ _1973_ VPWR VGND _1939_ sg13g2_nand4_1
X_4129_ _0968_ _0944_ _0967_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_58 VPWR VGND sg13g2_fill_1
XFILLER_40_845 VPWR VGND sg13g2_fill_1
XFILLER_8_518 VPWR VGND sg13g2_fill_2
XFILLER_40_878 VPWR VGND sg13g2_decap_8
XFILLER_4_779 VPWR VGND sg13g2_fill_1
Xfanout1002 DP_3.matrix\[8\] net1002 VPWR VGND sg13g2_buf_1
XFILLER_0_941 VPWR VGND sg13g2_decap_8
Xfanout1013 net1016 net1013 VPWR VGND sg13g2_buf_8
XFILLER_48_912 VPWR VGND sg13g2_decap_8
Xfanout1024 net1025 net1024 VPWR VGND sg13g2_buf_8
Xfanout1046 net1047 net1046 VPWR VGND sg13g2_buf_8
Xfanout1035 net1037 net1035 VPWR VGND sg13g2_buf_8
Xfanout1068 net1069 net1068 VPWR VGND sg13g2_buf_8
Xfanout1079 net1087 net1079 VPWR VGND sg13g2_buf_8
Xfanout1057 net1058 net1057 VPWR VGND sg13g2_buf_8
XFILLER_48_989 VPWR VGND sg13g2_decap_8
XFILLER_16_853 VPWR VGND sg13g2_fill_2
XFILLER_43_650 VPWR VGND sg13g2_fill_1
XFILLER_37_1014 VPWR VGND sg13g2_decap_8
XFILLER_31_878 VPWR VGND sg13g2_decap_8
X_3500_ _0362_ net931 net984 VPWR VGND sg13g2_nand2_1
X_4480_ _1304_ net803 net856 VPWR VGND sg13g2_nand2_1
Xhold507 _2114_ VPWR VGND net547 sg13g2_dlygate4sd3_1
X_3431_ _0295_ net931 net988 VPWR VGND sg13g2_nand2_1
X_3362_ _2948_ _2924_ _2947_ VPWR VGND sg13g2_xnor2_1
X_6150_ net1074 VGND VPWR _0255_ DP_4.matrix\[39\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_5101_ _1896_ _1897_ _1898_ VPWR VGND sg13g2_and2_1
X_6081_ net1079 VGND VPWR _0207_ DP_2.matrix\[39\] clknet_leaf_51_clk sg13g2_dfrbpq_2
X_3293_ _0096_ _2880_ _2881_ VPWR VGND sg13g2_xnor2_1
X_5032_ _1830_ _1825_ _1829_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_923 VPWR VGND sg13g2_decap_8
XFILLER_18_0 VPWR VGND sg13g2_fill_2
X_5934_ net951 _0192_ VPWR VGND sg13g2_buf_1
XFILLER_34_650 VPWR VGND sg13g2_fill_2
X_5865_ _2438_ _2436_ _2556_ VPWR VGND sg13g2_xor2_1
X_4816_ _1615_ _1625_ _1626_ VPWR VGND sg13g2_nor2_1
X_5796_ net829 _2463_ _2502_ VPWR VGND sg13g2_nor2_1
X_4747_ _1559_ _1544_ _1558_ VPWR VGND sg13g2_nand2_1
X_4678_ _1490_ _1451_ _1491_ VPWR VGND sg13g2_xor2_1
X_6417_ net1094 VGND VPWR net121 mac2.sum_lvl1_ff\[50\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3629_ _0488_ DP_2.matrix\[3\] net980 VPWR VGND sg13g2_nand2_1
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
X_6348_ net1091 VGND VPWR _0148_ mac2.products_ff\[9\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_6279_ net1022 VGND VPWR net142 mac1.sum_lvl3_ff\[24\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_45_937 VPWR VGND sg13g2_decap_8
XFILLER_44_447 VPWR VGND sg13g2_fill_2
XFILLER_16_149 VPWR VGND sg13g2_fill_1
XFILLER_25_650 VPWR VGND sg13g2_fill_1
XFILLER_31_119 VPWR VGND sg13g2_fill_1
XFILLER_9_805 VPWR VGND sg13g2_fill_2
XFILLER_9_838 VPWR VGND sg13g2_fill_2
XFILLER_8_304 VPWR VGND sg13g2_fill_2
XFILLER_4_521 VPWR VGND sg13g2_fill_1
XFILLER_48_764 VPWR VGND sg13g2_decap_8
XFILLER_35_425 VPWR VGND sg13g2_fill_2
XFILLER_36_948 VPWR VGND sg13g2_decap_8
XFILLER_44_970 VPWR VGND sg13g2_decap_8
X_3980_ _0823_ _0816_ _0824_ VPWR VGND sg13g2_xor2_1
X_5650_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] _2359_ VPWR VGND sg13g2_and2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_4601_ _1416_ _1408_ _1412_ VPWR VGND sg13g2_nand2_1
XFILLER_31_697 VPWR VGND sg13g2_fill_1
X_5581_ mac1.total_sum\[1\] mac2.total_sum\[1\] _2306_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_4532_ net833 net884 net829 net882 _1351_ VPWR VGND sg13g2_and4_1
Xhold304 DP_4.matrix\[4\] VPWR VGND net344 sg13g2_dlygate4sd3_1
X_4463_ _1287_ _1286_ _1288_ VPWR VGND sg13g2_nor2b_1
Xhold315 _0026_ VPWR VGND net355 sg13g2_dlygate4sd3_1
Xhold326 DP_4.matrix\[2\] VPWR VGND net366 sg13g2_dlygate4sd3_1
X_6202_ net1078 VGND VPWR net173 mac1.sum_lvl2_ff\[26\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3414_ _0277_ _0278_ _0272_ _0279_ VPWR VGND sg13g2_nand3_1
Xhold348 DP_2.matrix\[2\] VPWR VGND net388 sg13g2_dlygate4sd3_1
Xhold337 mac1.sum_lvl3_ff\[10\] VPWR VGND net377 sg13g2_dlygate4sd3_1
Xhold359 _2295_ VPWR VGND net399 sg13g2_dlygate4sd3_1
Xfanout806 net482 net806 VPWR VGND sg13g2_buf_8
X_4394_ net810 net807 net859 net856 _1221_ VPWR VGND sg13g2_and4_1
Xfanout839 net840 net839 VPWR VGND sg13g2_buf_1
Xfanout828 DP_4.matrix\[2\] net828 VPWR VGND sg13g2_buf_1
X_3345_ _2929_ _2912_ _2932_ VPWR VGND sg13g2_xor2_1
X_6133_ net1082 VGND VPWR net150 mac1.sum_lvl1_ff\[12\] clknet_leaf_43_clk sg13g2_dfrbpq_1
Xfanout817 net818 net817 VPWR VGND sg13g2_buf_2
X_6064_ net1014 VGND VPWR _0094_ mac1.products_ff\[141\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3276_ _2865_ net948 net887 VPWR VGND sg13g2_nand2_1
X_5015_ _1812_ _1784_ _1814_ VPWR VGND sg13g2_xor2_1
XFILLER_27_959 VPWR VGND sg13g2_decap_8
X_5917_ net275 _0165_ VPWR VGND sg13g2_buf_1
XFILLER_22_620 VPWR VGND sg13g2_fill_2
XFILLER_35_992 VPWR VGND sg13g2_decap_8
XFILLER_21_130 VPWR VGND sg13g2_fill_2
XFILLER_22_642 VPWR VGND sg13g2_fill_1
XFILLER_34_480 VPWR VGND sg13g2_fill_1
X_5848_ net932 net754 _2544_ VPWR VGND sg13g2_nor2_1
XFILLER_22_686 VPWR VGND sg13g2_decap_4
X_5779_ _2486_ _2483_ _2485_ VPWR VGND sg13g2_nand2b_1
XFILLER_10_859 VPWR VGND sg13g2_fill_1
XFILLER_10_848 VPWR VGND sg13g2_fill_1
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_29_274 VPWR VGND sg13g2_fill_2
XFILLER_26_992 VPWR VGND sg13g2_decap_8
XFILLER_41_962 VPWR VGND sg13g2_decap_8
XFILLER_34_1017 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_450 VPWR VGND sg13g2_fill_2
X_3130_ _2701_ _2720_ _2722_ _2723_ VPWR VGND sg13g2_or3_1
X_3061_ VGND VPWR _2654_ _2655_ _2656_ _2618_ sg13g2_a21oi_1
XFILLER_36_701 VPWR VGND sg13g2_decap_4
XFILLER_35_222 VPWR VGND sg13g2_fill_1
XFILLER_36_745 VPWR VGND sg13g2_fill_1
XFILLER_24_918 VPWR VGND sg13g2_fill_1
XFILLER_36_767 VPWR VGND sg13g2_decap_4
X_3963_ _0807_ _0800_ _0806_ VPWR VGND sg13g2_xnor2_1
X_3894_ _0740_ _0722_ _0738_ _0739_ VPWR VGND sg13g2_and3_1
X_5702_ VGND VPWR _2591_ net773 _2410_ _2409_ sg13g2_a21oi_1
XFILLER_32_962 VPWR VGND sg13g2_decap_8
X_5633_ _2347_ mac1.total_sum\[12\] mac2.total_sum\[12\] VPWR VGND sg13g2_nand2_1
X_5564_ net312 VPWR _2294_ VGND _2289_ _2290_ sg13g2_o21ai_1
X_4515_ _1324_ _1337_ _1338_ VPWR VGND sg13g2_nor2_1
Xhold101 mac2.sum_lvl1_ff\[48\] VPWR VGND net141 sg13g2_dlygate4sd3_1
Xhold134 mac2.sum_lvl2_ff\[53\] VPWR VGND net174 sg13g2_dlygate4sd3_1
X_5495_ _2240_ mac2.sum_lvl2_ff\[32\] mac2.sum_lvl2_ff\[13\] VPWR VGND sg13g2_xnor2_1
Xhold112 mac1.products_ff\[75\] VPWR VGND net152 sg13g2_dlygate4sd3_1
Xhold123 mac2.products_ff\[68\] VPWR VGND net163 sg13g2_dlygate4sd3_1
X_4446_ _1271_ net805 net1000 VPWR VGND sg13g2_nand2_2
Xhold167 mac1.sum_lvl1_ff\[82\] VPWR VGND net207 sg13g2_dlygate4sd3_1
Xhold145 mac2.products_ff\[141\] VPWR VGND net185 sg13g2_dlygate4sd3_1
Xhold156 mac2.sum_lvl1_ff\[72\] VPWR VGND net196 sg13g2_dlygate4sd3_1
Xhold178 mac2.products_ff\[74\] VPWR VGND net218 sg13g2_dlygate4sd3_1
Xhold189 mac2.products_ff\[73\] VPWR VGND net229 sg13g2_dlygate4sd3_1
X_4377_ _1173_ _1167_ _1175_ _1204_ VPWR VGND sg13g2_a21o_1
X_3328_ _2915_ net948 net1003 VPWR VGND sg13g2_nand2_1
X_6116_ net1074 VGND VPWR _0230_ DP_3.matrix\[38\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6047_ net1086 VGND VPWR _0184_ DP_1.matrix\[40\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_3259_ _2847_ _2848_ _2849_ VPWR VGND sg13g2_nor2b_1
XFILLER_42_726 VPWR VGND sg13g2_fill_2
XFILLER_41_214 VPWR VGND sg13g2_fill_1
XFILLER_26_299 VPWR VGND sg13g2_fill_2
XFILLER_23_984 VPWR VGND sg13g2_decap_8
XFILLER_2_800 VPWR VGND sg13g2_fill_1
XFILLER_1_310 VPWR VGND sg13g2_fill_2
XFILLER_45_542 VPWR VGND sg13g2_fill_2
XFILLER_17_222 VPWR VGND sg13g2_fill_2
XFILLER_33_715 VPWR VGND sg13g2_fill_1
XFILLER_33_737 VPWR VGND sg13g2_fill_2
XFILLER_41_781 VPWR VGND sg13g2_fill_1
X_5280_ _2070_ _2060_ _2071_ VPWR VGND sg13g2_nor2b_1
X_4300_ _1129_ _1085_ _1128_ VPWR VGND sg13g2_xnor2_1
X_4231_ _1062_ net812 net864 VPWR VGND sg13g2_nand2_1
X_4162_ _0991_ VPWR _0996_ VGND _0992_ _0994_ sg13g2_o21ai_1
XFILLER_49_870 VPWR VGND sg13g2_decap_8
X_3113_ _2706_ _2669_ _2704_ VPWR VGND sg13g2_xnor2_1
X_4093_ _0914_ _0907_ _0916_ _0933_ VPWR VGND sg13g2_a21o_1
X_3044_ _2638_ _2617_ _2639_ VPWR VGND sg13g2_xor2_1
XFILLER_36_597 VPWR VGND sg13g2_fill_2
X_4995_ _1794_ _1793_ _1790_ VPWR VGND sg13g2_nand2b_1
X_3946_ _0788_ _0789_ _0720_ _0791_ VPWR VGND sg13g2_nand3_1
X_3877_ _0723_ net973 net911 VPWR VGND sg13g2_nand2_1
X_5616_ mac1.total_sum\[9\] mac2.total_sum\[9\] _2333_ VPWR VGND sg13g2_nor2_1
XFILLER_20_998 VPWR VGND sg13g2_decap_8
X_5547_ _0063_ _2277_ net339 VPWR VGND sg13g2_xnor2_1
XFILLER_2_107 VPWR VGND sg13g2_fill_1
X_5478_ net544 mac2.sum_lvl2_ff\[29\] _2226_ VPWR VGND sg13g2_xor2_1
X_4429_ _1255_ _1209_ _1253_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_58 VPWR VGND sg13g2_fill_1
XFILLER_24_1016 VPWR VGND sg13g2_decap_8
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_328 VPWR VGND sg13g2_fill_1
XFILLER_7_936 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_49_133 VPWR VGND sg13g2_decap_8
XFILLER_18_597 VPWR VGND sg13g2_decap_8
X_4780_ _1586_ VPWR _1591_ VGND _1588_ _1589_ sg13g2_o21ai_1
X_3800_ _0649_ _0647_ _0648_ VPWR VGND sg13g2_nand2_1
XFILLER_33_567 VPWR VGND sg13g2_fill_1
X_3731_ _0109_ _0585_ _0586_ VPWR VGND sg13g2_xnor2_1
X_3662_ _0520_ net984 net926 VPWR VGND sg13g2_nand2_1
X_6450_ net1089 VGND VPWR net73 mac2.sum_lvl2_ff\[29\] clknet_leaf_37_clk sg13g2_dfrbpq_1
Xclkload10 clknet_4_13_0_clk clkload10/X VPWR VGND sg13g2_buf_8
X_5401_ net407 _2166_ _0030_ VPWR VGND sg13g2_nor2b_1
Xclkload21 VPWR clkload21/Y clknet_leaf_50_clk VGND sg13g2_inv_1
X_3593_ net934 net930 net979 net1010 _0453_ VPWR VGND sg13g2_and4_1
X_6381_ net1026 VGND VPWR _0150_ mac2.products_ff\[146\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5332_ mac1.sum_lvl2_ff\[28\] mac1.sum_lvl2_ff\[9\] _2113_ VPWR VGND sg13g2_nor2_1
XFILLER_47_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_1016 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_fill_2
X_5263_ _2053_ _2054_ _2055_ VPWR VGND sg13g2_nor2b_1
X_5194_ _1988_ net848 net994 VPWR VGND sg13g2_nand2_1
X_4214_ _1019_ _1043_ _1044_ _1046_ VPWR VGND sg13g2_nor3_1
X_4145_ _0981_ net869 net813 _0079_ VPWR VGND sg13g2_and3_2
X_4076_ _0915_ _0906_ _0917_ VPWR VGND sg13g2_xor2_1
X_3027_ net898 net952 net903 _2623_ VPWR VGND net949 sg13g2_nand4_1
XFILLER_37_895 VPWR VGND sg13g2_decap_8
XFILLER_24_578 VPWR VGND sg13g2_fill_2
X_4978_ VGND VPWR _1776_ _1777_ _1778_ _1740_ sg13g2_a21oi_1
X_3929_ net919 net960 net922 _0774_ VPWR VGND net1008 sg13g2_nand4_1
Xclkload4 clknet_4_6_0_clk clkload4/X VPWR VGND sg13g2_buf_8
XFILLER_3_449 VPWR VGND sg13g2_fill_1
XFILLER_28_895 VPWR VGND sg13g2_decap_8
XFILLER_24_82 VPWR VGND sg13g2_fill_2
XFILLER_40_81 VPWR VGND sg13g2_fill_2
XFILLER_49_90 VPWR VGND sg13g2_decap_8
XFILLER_38_604 VPWR VGND sg13g2_decap_4
X_5950_ net893 _0216_ VPWR VGND sg13g2_buf_1
X_4901_ _1707_ _1691_ _0143_ VPWR VGND sg13g2_xor2_1
XFILLER_19_895 VPWR VGND sg13g2_fill_1
X_5881_ _2476_ _2472_ _2566_ VPWR VGND sg13g2_xor2_1
X_4832_ _1612_ VPWR _1641_ VGND _1610_ _1613_ sg13g2_o21ai_1
XFILLER_33_375 VPWR VGND sg13g2_fill_2
XFILLER_34_898 VPWR VGND sg13g2_decap_8
X_4763_ _1547_ VPWR _1574_ VGND _1545_ _1548_ sg13g2_o21ai_1
X_3714_ _0570_ DP_2.matrix\[6\] net980 VPWR VGND sg13g2_nand2_1
X_4694_ net835 net832 net873 net1001 _1507_ VPWR VGND sg13g2_and4_1
X_6433_ net1090 VGND VPWR net200 mac2.sum_lvl2_ff\[9\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_3645_ VGND VPWR _0426_ _0467_ _0504_ _0468_ sg13g2_a21oi_1
X_3576_ _0436_ net988 net926 VPWR VGND sg13g2_nand2_1
X_6364_ net1088 VGND VPWR _0137_ mac2.products_ff\[77\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5315_ _0011_ _2097_ net530 VPWR VGND sg13g2_xnor2_1
X_6295_ net1023 VGND VPWR _0010_ mac1.sum_lvl3_ff\[4\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_5246_ _2038_ net844 net994 VPWR VGND sg13g2_nand2_1
XFILLER_29_27 VPWR VGND sg13g2_fill_2
Xhold16 mac2.sum_lvl2_ff\[49\] VPWR VGND net56 sg13g2_dlygate4sd3_1
Xhold38 mac2.products_ff\[3\] VPWR VGND net78 sg13g2_dlygate4sd3_1
Xhold27 mac2.sum_lvl2_ff\[45\] VPWR VGND net67 sg13g2_dlygate4sd3_1
Xhold49 mac1.products_ff\[0\] VPWR VGND net89 sg13g2_dlygate4sd3_1
X_5177_ _1970_ _1971_ _1972_ VPWR VGND sg13g2_nor2b_1
X_4128_ _0965_ _0964_ _0967_ VPWR VGND sg13g2_xor2_1
X_4059_ _0118_ _0899_ _0900_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_128 VPWR VGND sg13g2_fill_1
XFILLER_25_821 VPWR VGND sg13g2_decap_8
XFILLER_3_202 VPWR VGND sg13g2_fill_1
XFILLER_3_224 VPWR VGND sg13g2_fill_2
XFILLER_0_920 VPWR VGND sg13g2_decap_8
Xfanout1003 DP_2.matrix\[80\] net1003 VPWR VGND sg13g2_buf_8
Xfanout1047 net1048 net1047 VPWR VGND sg13g2_buf_8
Xfanout1014 net1016 net1014 VPWR VGND sg13g2_buf_8
Xfanout1025 net1098 net1025 VPWR VGND sg13g2_buf_8
Xfanout1036 net1037 net1036 VPWR VGND sg13g2_buf_8
XFILLER_0_997 VPWR VGND sg13g2_decap_8
Xfanout1069 net1071 net1069 VPWR VGND sg13g2_buf_8
Xfanout1058 net1059 net1058 VPWR VGND sg13g2_buf_8
XFILLER_48_968 VPWR VGND sg13g2_decap_8
XFILLER_47_445 VPWR VGND sg13g2_fill_1
XFILLER_35_607 VPWR VGND sg13g2_fill_1
XFILLER_7_530 VPWR VGND sg13g2_fill_2
Xhold508 mac1.sum_lvl2_ff\[10\] VPWR VGND net548 sg13g2_dlygate4sd3_1
X_3430_ _0275_ VPWR _0294_ VGND _0273_ _0276_ sg13g2_o21ai_1
X_3361_ _2945_ _2944_ _2947_ VPWR VGND sg13g2_xor2_1
XFILLER_44_1019 VPWR VGND sg13g2_decap_8
X_6080_ net1086 VGND VPWR _0206_ DP_2.matrix\[38\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_5100_ _1894_ _1893_ _1895_ _1897_ VPWR VGND sg13g2_a21o_1
X_3292_ VGND VPWR _2849_ _2852_ _2881_ _2847_ sg13g2_a21oi_1
XFILLER_39_902 VPWR VGND sg13g2_decap_8
X_5031_ _1829_ _1791_ _1827_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_423 VPWR VGND sg13g2_fill_2
XFILLER_39_979 VPWR VGND sg13g2_decap_8
X_5933_ net953 _0191_ VPWR VGND sg13g2_buf_1
XFILLER_15_29 VPWR VGND sg13g2_fill_1
X_5864_ net926 net755 _2555_ VPWR VGND sg13g2_nor2_1
XFILLER_21_301 VPWR VGND sg13g2_fill_2
X_4815_ _1623_ _1616_ _1625_ VPWR VGND sg13g2_xor2_1
X_5795_ _2501_ _2500_ net767 net765 net800 VPWR VGND sg13g2_a22oi_1
X_4746_ _1557_ _1550_ _1558_ VPWR VGND sg13g2_xor2_1
X_4677_ _1490_ net883 net821 VPWR VGND sg13g2_nand2_1
X_3628_ _0487_ DP_2.matrix\[4\] net980 VPWR VGND sg13g2_nand2_2
X_6416_ net1094 VGND VPWR net165 mac2.sum_lvl1_ff\[49\] clknet_leaf_36_clk sg13g2_dfrbpq_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
Xoutput17 net17 uio_out[0] VPWR VGND sg13g2_buf_1
X_6347_ net1088 VGND VPWR _0147_ mac2.products_ff\[8\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_3559_ _0395_ VPWR _0420_ VGND _0416_ _0418_ sg13g2_o21ai_1
X_6278_ net1039 VGND VPWR net260 mac1.sum_lvl3_ff\[23\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5229_ VGND VPWR _2022_ _2021_ _2010_ sg13g2_or2_1
XFILLER_45_916 VPWR VGND sg13g2_decap_8
XFILLER_31_109 VPWR VGND sg13g2_fill_1
XFILLER_13_846 VPWR VGND sg13g2_fill_2
XFILLER_4_511 VPWR VGND sg13g2_fill_1
XFILLER_36_927 VPWR VGND sg13g2_decap_8
X_4600_ _0138_ _1388_ _1415_ VPWR VGND sg13g2_xnor2_1
X_5580_ _2305_ mac1.total_sum\[1\] mac2.total_sum\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_7_63 VPWR VGND sg13g2_fill_1
X_4531_ net886 net827 _1350_ VPWR VGND sg13g2_and2_1
Xhold316 DP_4.matrix\[77\] VPWR VGND net356 sg13g2_dlygate4sd3_1
X_4462_ VGND VPWR _1242_ _1247_ _1287_ _1260_ sg13g2_a21oi_1
Xhold305 DP_2.matrix\[73\] VPWR VGND net345 sg13g2_dlygate4sd3_1
XFILLER_8_894 VPWR VGND sg13g2_fill_2
Xhold327 mac2.sum_lvl3_ff\[15\] VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold349 _0198_ VPWR VGND net389 sg13g2_dlygate4sd3_1
X_3413_ _0273_ VPWR _0278_ VGND _0274_ _0276_ sg13g2_o21ai_1
X_6201_ net1078 VGND VPWR net183 mac1.sum_lvl2_ff\[25\] clknet_leaf_51_clk sg13g2_dfrbpq_1
Xhold338 _2173_ VPWR VGND net378 sg13g2_dlygate4sd3_1
X_4393_ _1220_ net807 net856 VPWR VGND sg13g2_nand2_1
Xfanout807 net808 net807 VPWR VGND sg13g2_buf_8
X_3344_ _2912_ _2929_ _2931_ VPWR VGND sg13g2_nor2_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
Xfanout829 net359 net829 VPWR VGND sg13g2_buf_8
Xfanout818 DP_4.matrix\[36\] net818 VPWR VGND sg13g2_buf_2
X_6132_ net1056 VGND VPWR _0241_ DP_3.matrix\[77\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3275_ _2864_ net953 net1003 VPWR VGND sg13g2_nand2_1
X_6063_ net1047 VGND VPWR _0195_ DP_1.matrix\[79\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5014_ _1813_ _1784_ _1812_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_938 VPWR VGND sg13g2_decap_8
X_5916_ net1004 _0164_ VPWR VGND sg13g2_buf_1
XFILLER_35_971 VPWR VGND sg13g2_decap_8
X_5847_ net754 net937 _0196_ VPWR VGND sg13g2_xor2_1
X_5778_ _2485_ _2484_ net768 net766 net840 VPWR VGND sg13g2_a22oi_1
X_4729_ _1541_ _1534_ _1540_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_905 VPWR VGND sg13g2_decap_4
XFILLER_26_971 VPWR VGND sg13g2_decap_8
XFILLER_32_418 VPWR VGND sg13g2_fill_2
XFILLER_32_429 VPWR VGND sg13g2_fill_2
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_13_665 VPWR VGND sg13g2_decap_4
XFILLER_8_168 VPWR VGND sg13g2_fill_1
XFILLER_5_886 VPWR VGND sg13g2_decap_4
X_3060_ _2653_ _2652_ _2635_ _2655_ VPWR VGND sg13g2_a21o_1
XFILLER_35_234 VPWR VGND sg13g2_fill_1
XFILLER_17_982 VPWR VGND sg13g2_decap_8
X_5701_ net771 VPWR _2409_ VGND DP_2.matrix\[44\] net773 sg13g2_o21ai_1
X_3962_ _0805_ _0801_ _0806_ VPWR VGND sg13g2_xor2_1
XFILLER_16_470 VPWR VGND sg13g2_fill_1
XFILLER_32_941 VPWR VGND sg13g2_decap_8
X_3893_ _0727_ VPWR _0739_ VGND _0735_ _0737_ sg13g2_o21ai_1
X_5632_ _2344_ _2345_ _2346_ VPWR VGND sg13g2_nor2_1
X_5563_ net311 mac2.sum_lvl3_ff\[32\] _2293_ VPWR VGND sg13g2_xor2_1
X_4514_ _1335_ _1325_ _1337_ VPWR VGND sg13g2_xor2_1
Xhold113 mac1.sum_lvl1_ff\[77\] VPWR VGND net153 sg13g2_dlygate4sd3_1
Xhold102 mac1.sum_lvl2_ff\[42\] VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold135 mac1.products_ff\[141\] VPWR VGND net175 sg13g2_dlygate4sd3_1
Xhold124 mac1.sum_lvl1_ff\[83\] VPWR VGND net164 sg13g2_dlygate4sd3_1
X_5494_ _0035_ _2236_ _2238_ VPWR VGND sg13g2_xnor2_1
X_4445_ _1270_ net1000 net807 net856 net805 VPWR VGND sg13g2_a22oi_1
Xhold157 mac1.sum_lvl1_ff\[36\] VPWR VGND net197 sg13g2_dlygate4sd3_1
Xhold146 mac2.products_ff\[76\] VPWR VGND net186 sg13g2_dlygate4sd3_1
Xhold168 mac2.products_ff\[143\] VPWR VGND net208 sg13g2_dlygate4sd3_1
X_4376_ _1203_ _1202_ _0137_ VPWR VGND sg13g2_xor2_1
Xhold179 mac2.products_ff\[149\] VPWR VGND net219 sg13g2_dlygate4sd3_1
X_6115_ net1069 VGND VPWR net147 mac1.sum_lvl1_ff\[6\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3327_ _2893_ VPWR _2914_ VGND _2865_ _2891_ sg13g2_o21ai_1
X_6046_ net1079 VGND VPWR _0183_ DP_1.matrix\[39\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_3258_ _2810_ _2846_ _2808_ _2848_ VPWR VGND sg13g2_nand3_1
XFILLER_39_540 VPWR VGND sg13g2_fill_2
X_3189_ VGND VPWR _2780_ _2748_ _2746_ sg13g2_or2_1
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
XFILLER_26_201 VPWR VGND sg13g2_fill_1
XFILLER_27_746 VPWR VGND sg13g2_fill_2
XFILLER_41_237 VPWR VGND sg13g2_fill_2
XFILLER_10_602 VPWR VGND sg13g2_decap_4
XFILLER_23_963 VPWR VGND sg13g2_decap_8
XFILLER_10_624 VPWR VGND sg13g2_fill_1
XFILLER_2_878 VPWR VGND sg13g2_fill_2
XFILLER_40_1011 VPWR VGND sg13g2_decap_8
XFILLER_14_985 VPWR VGND sg13g2_decap_8
XFILLER_9_488 VPWR VGND sg13g2_decap_8
X_4230_ _1032_ VPWR _1061_ VGND _1030_ _1033_ sg13g2_o21ai_1
X_4161_ _0991_ _0992_ _0994_ _0995_ VPWR VGND sg13g2_nor3_1
X_3112_ VGND VPWR _2705_ _2704_ _2669_ sg13g2_or2_1
X_4092_ _0922_ _0901_ _0921_ _0932_ VPWR VGND sg13g2_a21o_1
X_3043_ _2638_ net954 net894 VPWR VGND sg13g2_nand2_1
XFILLER_36_576 VPWR VGND sg13g2_fill_2
XFILLER_23_215 VPWR VGND sg13g2_fill_1
X_4994_ _1792_ _1759_ _1793_ VPWR VGND sg13g2_xor2_1
X_3945_ _0789_ _0788_ _0720_ _0790_ VPWR VGND sg13g2_a21o_1
XFILLER_17_1024 VPWR VGND sg13g2_decap_4
X_3876_ _0703_ _0693_ _0701_ _0722_ VPWR VGND sg13g2_a21o_1
X_5615_ VGND VPWR mac1.total_sum\[8\] mac2.total_sum\[8\] _2332_ _2330_ sg13g2_a21oi_1
XFILLER_20_977 VPWR VGND sg13g2_decap_8
X_5546_ net338 mac2.sum_lvl3_ff\[29\] _2279_ VPWR VGND sg13g2_xor2_1
X_5477_ mac2.sum_lvl2_ff\[29\] mac2.sum_lvl2_ff\[10\] _2225_ VPWR VGND sg13g2_and2_1
X_4428_ VGND VPWR _1254_ _1252_ _1210_ sg13g2_or2_1
X_4359_ _1187_ net999 net815 net855 net811 VPWR VGND sg13g2_a22oi_1
X_6029_ net1075 VGND VPWR _0166_ DP_3.matrix\[8\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_42_513 VPWR VGND sg13g2_fill_1
XFILLER_42_579 VPWR VGND sg13g2_decap_8
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_13_62 VPWR VGND sg13g2_fill_2
XFILLER_49_156 VPWR VGND sg13g2_decap_8
Xfanout990 DP_1.matrix\[2\] net990 VPWR VGND sg13g2_buf_1
XFILLER_38_81 VPWR VGND sg13g2_fill_1
XFILLER_46_896 VPWR VGND sg13g2_decap_8
XFILLER_33_513 VPWR VGND sg13g2_fill_1
XFILLER_21_719 VPWR VGND sg13g2_fill_2
X_3730_ VGND VPWR _0560_ _0564_ _0586_ _0559_ sg13g2_a21oi_1
X_3661_ _0519_ net984 net925 VPWR VGND sg13g2_nand2_1
X_5400_ _2162_ net406 _2160_ _2166_ VPWR VGND sg13g2_nand3_1
X_3592_ _0452_ net931 net1010 VPWR VGND sg13g2_nand2_1
Xclkload11 clknet_4_14_0_clk clkload11/X VPWR VGND sg13g2_buf_8
X_6380_ net1027 VGND VPWR _0159_ mac2.products_ff\[145\] clknet_leaf_20_clk sg13g2_dfrbpq_1
Xclkload22 clkload22/Y clknet_leaf_31_clk VPWR VGND sg13g2_inv_2
X_5331_ VGND VPWR mac1.sum_lvl2_ff\[27\] mac1.sum_lvl2_ff\[8\] _2112_ _2110_ sg13g2_a21oi_1
X_5262_ _2054_ _2052_ _2035_ VPWR VGND sg13g2_nand2b_1
X_5193_ _1959_ VPWR _1987_ VGND _1956_ _1960_ sg13g2_o21ai_1
X_4213_ _1041_ _1042_ _1005_ _1045_ VPWR VGND sg13g2_nand3_1
X_4144_ net871 net819 _0079_ VPWR VGND sg13g2_and2_1
X_4075_ _0915_ _0906_ _0916_ VPWR VGND sg13g2_nor2b_1
X_3026_ net903 net899 net952 net949 _2622_ VPWR VGND sg13g2_and4_1
XFILLER_37_874 VPWR VGND sg13g2_decap_8
X_4977_ _1775_ _1774_ _1757_ _1777_ VPWR VGND sg13g2_a21o_1
X_3928_ net922 net919 net960 net1008 _0773_ VPWR VGND sg13g2_and4_1
Xclkload5 clknet_4_7_0_clk clkload5/X VPWR VGND sg13g2_buf_8
X_3859_ _0704_ _0705_ _0687_ _0706_ VPWR VGND sg13g2_nand3_1
X_5529_ mac2.sum_lvl3_ff\[26\] mac2.sum_lvl3_ff\[6\] _2265_ VPWR VGND sg13g2_and2_1
XFILLER_8_1022 VPWR VGND sg13g2_decap_8
XFILLER_47_638 VPWR VGND sg13g2_decap_4
XFILLER_43_811 VPWR VGND sg13g2_fill_2
XFILLER_28_874 VPWR VGND sg13g2_decap_8
XFILLER_42_321 VPWR VGND sg13g2_fill_2
XFILLER_43_899 VPWR VGND sg13g2_decap_8
XFILLER_10_240 VPWR VGND sg13g2_fill_1
XFILLER_7_745 VPWR VGND sg13g2_fill_1
XFILLER_6_233 VPWR VGND sg13g2_fill_2
XFILLER_6_277 VPWR VGND sg13g2_fill_1
XFILLER_41_8 VPWR VGND sg13g2_decap_4
XFILLER_3_984 VPWR VGND sg13g2_decap_8
X_4900_ _1705_ _1692_ _1707_ VPWR VGND sg13g2_xor2_1
X_5880_ _2565_ net878 net759 VPWR VGND sg13g2_nand2_1
X_4831_ _1620_ VPWR _1640_ VGND _1618_ _1621_ sg13g2_o21ai_1
XFILLER_33_354 VPWR VGND sg13g2_fill_2
XFILLER_34_877 VPWR VGND sg13g2_decap_8
XFILLER_21_538 VPWR VGND sg13g2_decap_4
X_4762_ _1538_ VPWR _1573_ VGND _1535_ _1539_ sg13g2_o21ai_1
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_3713_ _0569_ net980 DP_2.matrix\[7\] VPWR VGND sg13g2_nand2_1
X_4693_ _1506_ net828 net875 VPWR VGND sg13g2_nand2_1
X_3644_ _0383_ _0428_ _0382_ _0503_ VPWR VGND _0469_ sg13g2_nand4_1
X_6432_ net1090 VGND VPWR net227 mac2.sum_lvl2_ff\[8\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3575_ _0435_ net988 net925 VPWR VGND sg13g2_nand2_1
X_6363_ net1088 VGND VPWR _0136_ mac2.products_ff\[76\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5314_ net529 mac1.sum_lvl2_ff\[24\] _2099_ VPWR VGND sg13g2_xor2_1
X_6294_ net1039 VGND VPWR net496 mac1.sum_lvl3_ff\[3\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_5245_ _2017_ VPWR _2037_ VGND _1989_ _2015_ sg13g2_o21ai_1
Xhold28 mac1.products_ff\[3\] VPWR VGND net68 sg13g2_dlygate4sd3_1
Xhold17 mac1.products_ff\[2\] VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold39 mac2.products_ff\[71\] VPWR VGND net79 sg13g2_dlygate4sd3_1
X_5176_ _1934_ _1969_ _1932_ _1971_ VPWR VGND sg13g2_nand3_1
X_4127_ _0966_ _0964_ _0965_ VPWR VGND sg13g2_nand2_1
XFILLER_28_126 VPWR VGND sg13g2_fill_1
X_4058_ VGND VPWR _0869_ _0872_ _0900_ _0867_ sg13g2_a21oi_1
X_3009_ net898 net954 net904 _2606_ VPWR VGND net952 sg13g2_nand4_1
Xclkbuf_leaf_63_clk clknet_4_2_0_clk clknet_leaf_63_clk VPWR VGND sg13g2_buf_8
XFILLER_36_181 VPWR VGND sg13g2_fill_2
Xfanout1004 net390 net1004 VPWR VGND sg13g2_buf_8
Xfanout1015 net1016 net1015 VPWR VGND sg13g2_buf_1
Xfanout1026 net1030 net1026 VPWR VGND sg13g2_buf_8
Xfanout1037 net1038 net1037 VPWR VGND sg13g2_buf_8
Xfanout1048 net1063 net1048 VPWR VGND sg13g2_buf_8
XFILLER_0_976 VPWR VGND sg13g2_decap_8
Xfanout1059 net1062 net1059 VPWR VGND sg13g2_buf_8
XFILLER_48_947 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_54_clk clknet_4_8_0_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
XFILLER_16_855 VPWR VGND sg13g2_fill_1
XFILLER_15_365 VPWR VGND sg13g2_fill_2
XFILLER_7_575 VPWR VGND sg13g2_fill_2
XFILLER_7_564 VPWR VGND sg13g2_fill_1
X_3360_ _2946_ _2944_ _2945_ VPWR VGND sg13g2_nand2_1
X_3291_ _2878_ _2879_ _2880_ VPWR VGND sg13g2_nor2b_1
X_5030_ VGND VPWR _1828_ _1826_ _1792_ sg13g2_or2_1
XFILLER_18_2 VPWR VGND sg13g2_fill_1
XFILLER_39_958 VPWR VGND sg13g2_decap_8
XFILLER_26_619 VPWR VGND sg13g2_fill_2
X_5932_ net276 _0190_ VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_45_clk clknet_4_11_0_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
XFILLER_34_652 VPWR VGND sg13g2_fill_1
X_5863_ VGND VPWR net755 _2554_ _0201_ _2553_ sg13g2_a21oi_1
X_4814_ _1623_ _1616_ _1624_ VPWR VGND sg13g2_nor2b_1
X_5794_ net819 net833 net780 _2500_ VPWR VGND sg13g2_mux2_1
X_4745_ _1557_ _1551_ _1555_ VPWR VGND sg13g2_xnor2_1
X_4676_ _1489_ net883 net820 VPWR VGND sg13g2_nand2_1
X_3627_ _0486_ net984 net927 VPWR VGND sg13g2_nand2_1
X_6415_ net1091 VGND VPWR net167 mac2.sum_lvl1_ff\[48\] clknet_leaf_36_clk sg13g2_dfrbpq_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
X_3558_ _0395_ _0416_ _0418_ _0419_ VPWR VGND sg13g2_or3_1
Xoutput18 net18 uio_out[1] VPWR VGND sg13g2_buf_1
X_6346_ net1076 VGND VPWR _0146_ mac2.products_ff\[7\] clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_0_228 VPWR VGND sg13g2_fill_1
X_6277_ net1041 VGND VPWR net171 mac1.sum_lvl3_ff\[22\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3489_ _0348_ _0350_ _0351_ VPWR VGND sg13g2_nor2b_1
X_5228_ _2019_ _2011_ _2021_ VPWR VGND sg13g2_xor2_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
X_5159_ _1926_ VPWR _1954_ VGND _1920_ _1927_ sg13g2_o21ai_1
XFILLER_29_424 VPWR VGND sg13g2_fill_2
XFILLER_38_991 VPWR VGND sg13g2_decap_8
XFILLER_44_449 VPWR VGND sg13g2_fill_1
XFILLER_37_490 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_36_clk clknet_4_15_0_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_12_335 VPWR VGND sg13g2_fill_2
XFILLER_40_644 VPWR VGND sg13g2_fill_1
XFILLER_8_328 VPWR VGND sg13g2_fill_1
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_36_906 VPWR VGND sg13g2_decap_8
XFILLER_35_427 VPWR VGND sg13g2_fill_1
XFILLER_16_652 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_27_clk clknet_4_7_0_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_43_493 VPWR VGND sg13g2_fill_2
XFILLER_30_143 VPWR VGND sg13g2_fill_2
XFILLER_31_677 VPWR VGND sg13g2_decap_4
XFILLER_30_176 VPWR VGND sg13g2_fill_2
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
X_4530_ _1348_ _1349_ _0085_ VPWR VGND sg13g2_nor2_1
X_4461_ _1284_ _1273_ _1286_ VPWR VGND sg13g2_xor2_1
Xhold317 DP_2.matrix\[77\] VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold306 DP_2.matrix\[79\] VPWR VGND net346 sg13g2_dlygate4sd3_1
X_3412_ _0273_ _0274_ _0276_ _0277_ VPWR VGND sg13g2_or3_1
X_6200_ net1078 VGND VPWR net41 mac1.sum_lvl2_ff\[24\] clknet_leaf_50_clk sg13g2_dfrbpq_2
Xhold339 _0017_ VPWR VGND net379 sg13g2_dlygate4sd3_1
Xhold328 _2303_ VPWR VGND net368 sg13g2_dlygate4sd3_1
X_4392_ _1219_ net861 net805 VPWR VGND sg13g2_nand2_1
X_6131_ net1055 VGND VPWR _0240_ DP_3.matrix\[76\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3343_ _2930_ _2912_ _2929_ VPWR VGND sg13g2_nand2_1
Xfanout819 net337 net819 VPWR VGND sg13g2_buf_8
Xfanout808 net314 net808 VPWR VGND sg13g2_buf_8
X_3274_ VGND VPWR _2863_ _2836_ _2834_ sg13g2_or2_1
X_6062_ net1046 VGND VPWR _0194_ DP_1.matrix\[78\] clknet_leaf_59_clk sg13g2_dfrbpq_2
X_5013_ _1812_ _1788_ _1811_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_38_254 VPWR VGND sg13g2_fill_2
XFILLER_39_766 VPWR VGND sg13g2_decap_8
XFILLER_38_276 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_18_clk clknet_4_4_0_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_35_950 VPWR VGND sg13g2_decap_8
X_5915_ net269 _0162_ VPWR VGND sg13g2_buf_1
XFILLER_22_611 VPWR VGND sg13g2_decap_4
X_5846_ _2542_ VPWR _0179_ VGND _2407_ _2543_ sg13g2_o21ai_1
XFILLER_22_622 VPWR VGND sg13g2_fill_1
X_5777_ net857 net873 _2448_ _2484_ VPWR VGND sg13g2_mux2_1
XFILLER_10_828 VPWR VGND sg13g2_fill_1
XFILLER_21_176 VPWR VGND sg13g2_decap_8
X_2989_ VPWR DP_1.Q_range.data_plus_4\[6\] net8 VGND sg13g2_inv_1
X_4728_ _1539_ _1535_ _1540_ VPWR VGND sg13g2_xor2_1
X_4659_ _1461_ VPWR _1473_ VGND _1469_ _1471_ sg13g2_o21ai_1
X_6329_ net1013 VGND VPWR net486 mac1.total_sum\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_29_276 VPWR VGND sg13g2_fill_1
XFILLER_45_758 VPWR VGND sg13g2_fill_2
XFILLER_26_950 VPWR VGND sg13g2_decap_8
XFILLER_33_909 VPWR VGND sg13g2_decap_8
XFILLER_41_920 VPWR VGND sg13g2_decap_8
XFILLER_40_452 VPWR VGND sg13g2_fill_1
XFILLER_41_997 VPWR VGND sg13g2_decap_8
X_3961_ _0805_ _0755_ _0803_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_961 VPWR VGND sg13g2_decap_8
X_5700_ VGND VPWR _2376_ _2407_ _0160_ _2408_ sg13g2_a21oi_1
XFILLER_32_920 VPWR VGND sg13g2_decap_8
X_3892_ _0727_ _0735_ _0737_ _0738_ VPWR VGND sg13g2_or3_1
X_5631_ _2340_ _2335_ _2339_ _2345_ VPWR VGND sg13g2_a21o_1
XFILLER_32_997 VPWR VGND sg13g2_decap_8
X_5562_ _2292_ mac2.sum_lvl3_ff\[32\] net311 VPWR VGND sg13g2_nand2_1
X_4513_ _1335_ _1325_ _1336_ VPWR VGND sg13g2_nor2b_1
Xhold125 mac2.products_ff\[81\] VPWR VGND net165 sg13g2_dlygate4sd3_1
Xhold103 mac1.sum_lvl2_ff\[45\] VPWR VGND net143 sg13g2_dlygate4sd3_1
Xhold114 mac2.sum_lvl1_ff\[83\] VPWR VGND net154 sg13g2_dlygate4sd3_1
X_5493_ _2238_ VPWR _2239_ VGND _2234_ _2235_ sg13g2_o21ai_1
X_4444_ _1256_ _1250_ _1258_ _1269_ VPWR VGND sg13g2_a21o_1
Xhold147 mac1.sum_lvl1_ff\[3\] VPWR VGND net187 sg13g2_dlygate4sd3_1
Xhold158 mac1.products_ff\[1\] VPWR VGND net198 sg13g2_dlygate4sd3_1
Xhold136 mac1.products_ff\[147\] VPWR VGND net176 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold169 mac2.products_ff\[147\] VPWR VGND net209 sg13g2_dlygate4sd3_1
X_4375_ _1203_ _1160_ _1163_ VPWR VGND sg13g2_nand2_1
X_3326_ _2894_ _2888_ _2896_ _2913_ VPWR VGND sg13g2_a21o_1
X_6114_ net1057 VGND VPWR _0229_ DP_3.matrix\[37\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6045_ net1079 VGND VPWR _0182_ DP_1.matrix\[38\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3257_ VGND VPWR _2808_ _2810_ _2847_ _2846_ sg13g2_a21oi_1
XFILLER_2_1006 VPWR VGND sg13g2_decap_8
X_3188_ _2738_ VPWR _2779_ VGND _2697_ _2736_ sg13g2_o21ai_1
X_5829_ _2390_ _2393_ _2389_ _2532_ VPWR VGND sg13g2_nand3_1
XFILLER_1_312 VPWR VGND sg13g2_fill_1
XFILLER_45_544 VPWR VGND sg13g2_fill_1
XFILLER_17_224 VPWR VGND sg13g2_fill_1
XFILLER_45_599 VPWR VGND sg13g2_fill_2
XFILLER_14_964 VPWR VGND sg13g2_decap_8
XFILLER_41_761 VPWR VGND sg13g2_fill_1
X_4160_ _0994_ net865 net819 net867 net813 VPWR VGND sg13g2_a22oi_1
X_3111_ _2704_ net894 net950 VPWR VGND sg13g2_nand2_1
X_4091_ _0930_ _0926_ _0119_ VPWR VGND sg13g2_xor2_1
X_3042_ _2637_ net955 net892 VPWR VGND sg13g2_nand2_1
XFILLER_36_500 VPWR VGND sg13g2_fill_2
X_4993_ _1792_ net848 net789 VPWR VGND sg13g2_nand2_1
X_3944_ _0787_ _0786_ _0752_ _0789_ VPWR VGND sg13g2_a21o_1
XFILLER_17_1003 VPWR VGND sg13g2_decap_8
X_3875_ _0721_ _0715_ _0719_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_923 VPWR VGND sg13g2_fill_2
X_5614_ _2330_ _2331_ net17 VPWR VGND sg13g2_nor2b_1
XFILLER_31_282 VPWR VGND sg13g2_fill_1
X_5545_ mac2.sum_lvl3_ff\[29\] net338 _2278_ VPWR VGND sg13g2_nor2_1
X_5476_ _0047_ _2222_ net543 VPWR VGND sg13g2_xnor2_1
X_4427_ _1253_ net861 net803 VPWR VGND sg13g2_nand2_1
X_4358_ net815 net811 net855 net999 _1186_ VPWR VGND sg13g2_and4_1
X_3309_ _2895_ _2887_ _2897_ VPWR VGND sg13g2_xor2_1
X_4289_ _1117_ _1116_ _0135_ VPWR VGND sg13g2_xor2_1
X_6028_ net1048 VGND VPWR _0165_ DP_2.matrix\[80\] clknet_leaf_60_clk sg13g2_dfrbpq_2
XFILLER_27_500 VPWR VGND sg13g2_fill_2
XFILLER_11_956 VPWR VGND sg13g2_decap_8
XFILLER_49_146 VPWR VGND sg13g2_decap_4
Xfanout991 net392 net991 VPWR VGND sg13g2_buf_8
Xfanout980 net505 net980 VPWR VGND sg13g2_buf_8
XFILLER_46_875 VPWR VGND sg13g2_decap_8
XFILLER_45_363 VPWR VGND sg13g2_fill_1
XFILLER_18_588 VPWR VGND sg13g2_fill_1
XFILLER_13_271 VPWR VGND sg13g2_fill_1
X_3660_ _0518_ net988 net1005 VPWR VGND sg13g2_nand2_1
Xclkload23 VPWR clkload23/Y clknet_leaf_33_clk VGND sg13g2_inv_1
X_3591_ _0407_ VPWR _0451_ VGND _0405_ _0408_ sg13g2_o21ai_1
Xclkload12 clknet_4_15_0_clk clkload12/X VPWR VGND sg13g2_buf_8
XFILLER_6_982 VPWR VGND sg13g2_decap_8
X_5330_ _2110_ _2111_ _0014_ VPWR VGND sg13g2_nor2b_2
X_5261_ _2052_ _2035_ _2053_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_2 VPWR VGND sg13g2_fill_1
X_4212_ _1044_ _1005_ _1041_ _1042_ VPWR VGND sg13g2_and3_1
X_5192_ VPWR _1986_ _1985_ VGND sg13g2_inv_1
X_4143_ _0122_ _0973_ _0980_ VPWR VGND sg13g2_xnor2_1
X_4074_ _0915_ _0907_ _0914_ VPWR VGND sg13g2_xnor2_1
X_3025_ _2621_ net954 net896 VPWR VGND sg13g2_nand2_1
XFILLER_24_536 VPWR VGND sg13g2_fill_2
XFILLER_12_709 VPWR VGND sg13g2_fill_2
X_4976_ _1774_ _1775_ _1757_ _1776_ VPWR VGND sg13g2_nand3_1
X_3927_ _0772_ net916 net963 VPWR VGND sg13g2_nand2_1
X_3858_ _0703_ _0702_ _0693_ _0705_ VPWR VGND sg13g2_a21o_1
Xclkload6 clknet_4_9_0_clk clkload6/X VPWR VGND sg13g2_buf_8
X_3789_ _0622_ _0637_ _0638_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1011 VPWR VGND sg13g2_decap_8
XFILLER_4_919 VPWR VGND sg13g2_decap_8
X_5528_ _0059_ _2262_ net419 VPWR VGND sg13g2_xnor2_1
X_5459_ _2211_ mac2.sum_lvl2_ff\[25\] net524 VPWR VGND sg13g2_xnor2_1
XFILLER_8_1001 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_fill_1
XFILLER_46_127 VPWR VGND sg13g2_fill_2
XFILLER_28_853 VPWR VGND sg13g2_decap_8
XFILLER_43_878 VPWR VGND sg13g2_decap_8
XFILLER_24_84 VPWR VGND sg13g2_fill_1
XFILLER_3_963 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_fill_1
XFILLER_46_650 VPWR VGND sg13g2_fill_1
XFILLER_18_330 VPWR VGND sg13g2_fill_2
XFILLER_45_171 VPWR VGND sg13g2_fill_2
X_4830_ _1639_ _1638_ _1636_ VPWR VGND sg13g2_nand2b_1
X_4761_ _1559_ VPWR _1572_ VGND _1543_ _1560_ sg13g2_o21ai_1
XFILLER_14_1006 VPWR VGND sg13g2_decap_8
X_3712_ _0568_ net984 net1005 VPWR VGND sg13g2_nand2_1
X_4692_ _1465_ VPWR _1505_ VGND _1463_ _1466_ sg13g2_o21ai_1
X_3643_ _0500_ _0501_ _0502_ VPWR VGND sg13g2_nor2b_1
X_6431_ net1088 VGND VPWR net105 mac2.sum_lvl2_ff\[7\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6362_ net1088 VGND VPWR _0135_ mac2.products_ff\[75\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5313_ mac1.sum_lvl2_ff\[24\] mac1.sum_lvl2_ff\[5\] _2098_ VPWR VGND sg13g2_nor2_1
X_3574_ _0434_ net992 net1005 VPWR VGND sg13g2_nand2_1
X_6293_ net1041 VGND VPWR net417 mac1.sum_lvl3_ff\[2\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_5244_ _2018_ _2012_ _2020_ _2036_ VPWR VGND sg13g2_a21o_1
Xhold18 mac1.sum_lvl2_ff\[47\] VPWR VGND net58 sg13g2_dlygate4sd3_1
Xhold29 mac2.sum_lvl1_ff\[40\] VPWR VGND net69 sg13g2_dlygate4sd3_1
XFILLER_29_29 VPWR VGND sg13g2_fill_1
X_5175_ VGND VPWR _1932_ _1934_ _1970_ _1969_ sg13g2_a21oi_1
X_4126_ _0939_ VPWR _0965_ VGND _0909_ _0937_ sg13g2_o21ai_1
X_4057_ _0897_ _0898_ _0899_ VPWR VGND sg13g2_nor2b_1
X_3008_ net903 net899 net954 net952 _2605_ VPWR VGND sg13g2_and4_1
XFILLER_12_528 VPWR VGND sg13g2_decap_4
XFILLER_25_889 VPWR VGND sg13g2_decap_8
X_4959_ _1759_ net850 net787 VPWR VGND sg13g2_nand2_1
XFILLER_3_226 VPWR VGND sg13g2_fill_1
XFILLER_0_955 VPWR VGND sg13g2_decap_8
Xfanout1016 net1025 net1016 VPWR VGND sg13g2_buf_8
Xfanout1005 net490 net1005 VPWR VGND sg13g2_buf_8
Xfanout1027 net1030 net1027 VPWR VGND sg13g2_buf_8
Xfanout1038 net1098 net1038 VPWR VGND sg13g2_buf_8
XFILLER_48_926 VPWR VGND sg13g2_decap_8
XFILLER_19_105 VPWR VGND sg13g2_fill_2
Xfanout1049 net1053 net1049 VPWR VGND sg13g2_buf_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_532 VPWR VGND sg13g2_fill_1
XFILLER_3_771 VPWR VGND sg13g2_fill_1
X_3290_ _2845_ _2877_ _2843_ _2879_ VPWR VGND sg13g2_nand3_1
XFILLER_39_937 VPWR VGND sg13g2_decap_8
XFILLER_38_425 VPWR VGND sg13g2_fill_1
XFILLER_26_609 VPWR VGND sg13g2_fill_1
XFILLER_47_981 VPWR VGND sg13g2_decap_8
X_5931_ net957 _0189_ VPWR VGND sg13g2_buf_1
X_5862_ _2435_ _2413_ _2554_ VPWR VGND sg13g2_xor2_1
XFILLER_21_303 VPWR VGND sg13g2_fill_1
X_4813_ _1623_ _1617_ _1622_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_185 VPWR VGND sg13g2_fill_1
X_5793_ _2499_ _2498_ net769 net765 net790 VPWR VGND sg13g2_a22oi_1
XFILLER_21_358 VPWR VGND sg13g2_fill_2
X_4744_ _1556_ _1551_ _1555_ VPWR VGND sg13g2_nand2_1
XFILLER_30_892 VPWR VGND sg13g2_decap_8
X_4675_ _1488_ DP_3.matrix\[0\] net996 VPWR VGND sg13g2_nand2_1
X_3626_ VGND VPWR net933 net978 _0485_ _0452_ sg13g2_a21oi_1
X_6414_ net1089 VGND VPWR net112 mac2.sum_lvl1_ff\[47\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_3557_ VGND VPWR _0414_ _0415_ _0418_ _0396_ sg13g2_a21oi_1
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
X_6345_ net1073 VGND VPWR _0145_ mac2.products_ff\[6\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6276_ net1041 VGND VPWR net70 mac1.sum_lvl3_ff\[21\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_5227_ _2019_ _2011_ _2020_ VPWR VGND sg13g2_nor2b_1
X_3488_ VGND VPWR _0350_ _0349_ _0316_ sg13g2_or2_1
X_5158_ _1951_ _1943_ _1953_ VPWR VGND sg13g2_xor2_1
X_4109_ _0947_ _0933_ _0949_ VPWR VGND sg13g2_xor2_1
X_5089_ _1886_ _1866_ _1884_ _1885_ VPWR VGND sg13g2_and3_1
XFILLER_38_970 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_778 VPWR VGND sg13g2_decap_8
XFILLER_44_984 VPWR VGND sg13g2_decap_8
X_4460_ VGND VPWR _1285_ _1284_ _1273_ sg13g2_or2_1
Xhold307 mac2.sum_lvl3_ff\[14\] VPWR VGND net347 sg13g2_dlygate4sd3_1
Xhold318 DP_1.matrix\[0\] VPWR VGND net358 sg13g2_dlygate4sd3_1
X_3411_ _0276_ net985 net939 net987 net936 VPWR VGND sg13g2_a22oi_1
Xhold329 _0054_ VPWR VGND net369 sg13g2_dlygate4sd3_1
X_4391_ VGND VPWR net815 net855 _1218_ _1185_ sg13g2_a21oi_1
X_3342_ _2927_ _2913_ _2929_ VPWR VGND sg13g2_xor2_1
X_6130_ net1080 VGND VPWR net99 mac1.sum_lvl1_ff\[11\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_3_590 VPWR VGND sg13g2_fill_2
XFILLER_30_2 VPWR VGND sg13g2_fill_1
Xfanout809 net328 net809 VPWR VGND sg13g2_buf_8
X_6061_ net1014 VGND VPWR _0068_ mac1.products_ff\[140\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3273_ _2824_ VPWR _2862_ VGND _2821_ _2825_ sg13g2_o21ai_1
X_5012_ _1811_ _1808_ _1810_ VPWR VGND sg13g2_nand2_1
XFILLER_16_0 VPWR VGND sg13g2_fill_1
X_5914_ net1009 _0161_ VPWR VGND sg13g2_buf_1
XFILLER_34_450 VPWR VGND sg13g2_fill_1
XFILLER_34_461 VPWR VGND sg13g2_decap_4
X_5845_ _2404_ _2406_ _2543_ VPWR VGND sg13g2_and2_1
XFILLER_34_494 VPWR VGND sg13g2_decap_4
X_5776_ _2478_ _2482_ _2483_ VPWR VGND sg13g2_nor2b_1
X_2988_ VPWR DP_3.Q_range.data_plus_4\[6\] net12 VGND sg13g2_inv_1
X_4727_ _1539_ _1489_ _1537_ VPWR VGND sg13g2_xnor2_1
X_4658_ _1461_ _1469_ _1471_ _1472_ VPWR VGND sg13g2_or3_1
X_3609_ _0466_ _0468_ _0469_ VPWR VGND sg13g2_nor2_1
X_4589_ VGND VPWR _1401_ _1402_ _1405_ _1396_ sg13g2_a21oi_1
X_6328_ net1012 VGND VPWR net319 mac1.total_sum\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_6259_ net1052 VGND VPWR net77 mac2.sum_lvl1_ff\[72\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_45_748 VPWR VGND sg13g2_fill_2
XFILLER_32_409 VPWR VGND sg13g2_fill_1
XFILLER_13_634 VPWR VGND sg13g2_fill_2
XFILLER_41_976 VPWR VGND sg13g2_decap_8
XFILLER_32_51 VPWR VGND sg13g2_fill_2
XFILLER_40_497 VPWR VGND sg13g2_decap_8
XFILLER_10_1020 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_fill_2
XFILLER_36_726 VPWR VGND sg13g2_fill_2
X_3960_ VGND VPWR _0804_ _0802_ _0756_ sg13g2_or2_1
X_3891_ VGND VPWR _0733_ _0734_ _0737_ _0728_ sg13g2_a21oi_1
XFILLER_32_976 VPWR VGND sg13g2_decap_8
X_5630_ _2333_ _2337_ _2343_ _2344_ VPWR VGND sg13g2_nor3_1
X_5561_ _2289_ _2290_ _2291_ VPWR VGND sg13g2_nor2_1
X_4512_ _1335_ _1311_ _1334_ VPWR VGND sg13g2_xnor2_1
X_5492_ mac2.sum_lvl2_ff\[12\] mac2.sum_lvl2_ff\[31\] _2238_ VPWR VGND sg13g2_xor2_1
Xhold126 mac1.products_ff\[143\] VPWR VGND net166 sg13g2_dlygate4sd3_1
Xhold104 mac1.products_ff\[142\] VPWR VGND net144 sg13g2_dlygate4sd3_1
Xhold115 mac2.sum_lvl1_ff\[38\] VPWR VGND net155 sg13g2_dlygate4sd3_1
Xhold159 mac2.products_ff\[151\] VPWR VGND net199 sg13g2_dlygate4sd3_1
Xhold137 mac1.products_ff\[73\] VPWR VGND net177 sg13g2_dlygate4sd3_1
Xhold148 mac2.sum_lvl1_ff\[39\] VPWR VGND net188 sg13g2_dlygate4sd3_1
X_4443_ _0129_ _1267_ _1268_ VPWR VGND sg13g2_xnor2_1
X_4374_ _1199_ _1201_ _1202_ VPWR VGND sg13g2_nor2_1
X_3325_ _2902_ _2882_ _2901_ _2912_ VPWR VGND sg13g2_a21o_1
X_6113_ net1057 VGND VPWR _0228_ DP_3.matrix\[36\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_6044_ net1079 VGND VPWR _0181_ DP_1.matrix\[37\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_3256_ _2846_ _2817_ _2844_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_542 VPWR VGND sg13g2_fill_1
X_3187_ _2764_ VPWR _2778_ VGND _2742_ _2765_ sg13g2_o21ai_1
XFILLER_39_564 VPWR VGND sg13g2_fill_2
XFILLER_26_247 VPWR VGND sg13g2_fill_2
XFILLER_35_770 VPWR VGND sg13g2_fill_1
XFILLER_41_239 VPWR VGND sg13g2_fill_1
X_5828_ net989 net753 _2531_ VPWR VGND sg13g2_nor2_1
XFILLER_23_998 VPWR VGND sg13g2_decap_8
XFILLER_10_637 VPWR VGND sg13g2_fill_2
X_5759_ net852 net767 _2466_ VPWR VGND sg13g2_nor2_1
XFILLER_33_707 VPWR VGND sg13g2_fill_1
XFILLER_14_943 VPWR VGND sg13g2_decap_8
XFILLER_40_261 VPWR VGND sg13g2_fill_2
XFILLER_43_94 VPWR VGND sg13g2_decap_4
X_3110_ _2703_ net955 net890 VPWR VGND sg13g2_nand2_1
X_4090_ _0931_ _0926_ _0930_ VPWR VGND sg13g2_nand2_1
XFILLER_49_884 VPWR VGND sg13g2_decap_8
X_3041_ _2636_ net958 net890 VPWR VGND sg13g2_nand2_1
XFILLER_48_383 VPWR VGND sg13g2_fill_1
XFILLER_17_792 VPWR VGND sg13g2_fill_2
X_4992_ _1791_ net848 net787 VPWR VGND sg13g2_nand2_1
X_3943_ _0786_ _0787_ _0752_ _0788_ VPWR VGND sg13g2_nand3_1
XFILLER_16_280 VPWR VGND sg13g2_fill_1
X_3874_ _0715_ _0719_ _0720_ VPWR VGND sg13g2_and2_1
X_5613_ _2327_ _2329_ _2325_ _2331_ VPWR VGND sg13g2_nand3_1
XFILLER_9_980 VPWR VGND sg13g2_decap_8
X_5544_ VGND VPWR mac2.sum_lvl3_ff\[28\] mac2.sum_lvl3_ff\[8\] _2277_ _2275_ sg13g2_a21oi_1
X_5475_ net542 mac2.sum_lvl2_ff\[28\] _2224_ VPWR VGND sg13g2_xor2_1
X_4426_ _1252_ net861 net802 VPWR VGND sg13g2_nand2_1
X_4357_ _1185_ net812 net999 VPWR VGND sg13g2_nand2_1
X_3308_ _2895_ _2887_ _2896_ VPWR VGND sg13g2_nor2b_1
X_4288_ _1118_ _1116_ _1117_ VPWR VGND sg13g2_nand2_1
X_3239_ _2827_ _2819_ _2829_ VPWR VGND sg13g2_xor2_1
X_6027_ net1080 VGND VPWR _0164_ DP_2.matrix\[44\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_39_383 VPWR VGND sg13g2_fill_1
Xhold490 _2099_ VPWR VGND net530 sg13g2_dlygate4sd3_1
XFILLER_2_655 VPWR VGND sg13g2_decap_4
Xfanout970 DP_1.matrix\[40\] net970 VPWR VGND sg13g2_buf_8
Xfanout992 DP_1.matrix\[1\] net992 VPWR VGND sg13g2_buf_1
Xfanout981 net982 net981 VPWR VGND sg13g2_buf_8
XFILLER_18_534 VPWR VGND sg13g2_fill_2
XFILLER_33_537 VPWR VGND sg13g2_fill_2
XFILLER_9_265 VPWR VGND sg13g2_fill_2
Xclkload13 VPWR clkload13/Y clknet_leaf_65_clk VGND sg13g2_inv_1
X_3590_ _0450_ _0444_ _0449_ VPWR VGND sg13g2_xnor2_1
Xclkload24 clkload24/Y clknet_leaf_38_clk VPWR VGND sg13g2_inv_8
XFILLER_6_961 VPWR VGND sg13g2_decap_8
X_5260_ _2052_ _2036_ _2050_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_471 VPWR VGND sg13g2_fill_2
X_4211_ VGND VPWR _1041_ _1042_ _1043_ _1005_ sg13g2_a21oi_1
X_5191_ _1948_ VPWR _1985_ VGND _1945_ _1949_ sg13g2_o21ai_1
X_4142_ _0980_ _0974_ _0979_ VPWR VGND sg13g2_xnor2_1
X_4073_ _0914_ _0908_ _0913_ VPWR VGND sg13g2_xnor2_1
X_3024_ _2606_ VPWR _2620_ VGND _2604_ _2607_ sg13g2_o21ai_1
X_4975_ _1763_ VPWR _1775_ VGND _1771_ _1773_ sg13g2_o21ai_1
X_3926_ _0731_ VPWR _0771_ VGND _0729_ _0732_ sg13g2_o21ai_1
XFILLER_11_209 VPWR VGND sg13g2_fill_1
X_3857_ _0702_ _0703_ _0693_ _0704_ VPWR VGND sg13g2_nand3_1
Xclkload7 clknet_4_10_0_clk clkload7/X VPWR VGND sg13g2_buf_8
X_3788_ _0637_ net975 net913 VPWR VGND sg13g2_nand2_2
X_5527_ net418 mac2.sum_lvl3_ff\[25\] _2264_ VPWR VGND sg13g2_xor2_1
X_5458_ mac2.sum_lvl2_ff\[25\] mac2.sum_lvl2_ff\[6\] _2210_ VPWR VGND sg13g2_and2_1
X_5389_ VPWR VGND _2151_ _2150_ _2149_ mac1.sum_lvl3_ff\[25\] _2157_ mac1.sum_lvl3_ff\[5\]
+ sg13g2_a221oi_1
X_4409_ _1234_ _1235_ _1236_ VPWR VGND sg13g2_nor2b_1
XFILLER_42_323 VPWR VGND sg13g2_fill_1
XFILLER_42_356 VPWR VGND sg13g2_fill_2
XFILLER_10_297 VPWR VGND sg13g2_fill_1
XFILLER_40_95 VPWR VGND sg13g2_fill_1
XFILLER_3_942 VPWR VGND sg13g2_decap_8
XFILLER_19_843 VPWR VGND sg13g2_fill_2
XFILLER_18_375 VPWR VGND sg13g2_fill_1
XFILLER_33_356 VPWR VGND sg13g2_fill_1
X_4760_ _1540_ _1534_ _1542_ _1571_ VPWR VGND sg13g2_a21o_1
X_3711_ _0547_ VPWR _0567_ VGND _0519_ _0545_ sg13g2_o21ai_1
X_4691_ _1504_ _1503_ _1502_ VPWR VGND sg13g2_nand2b_1
X_3642_ _0464_ _0499_ _0462_ _0501_ VPWR VGND sg13g2_nand3_1
X_6430_ net1071 VGND VPWR net108 mac2.sum_lvl2_ff\[6\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_6361_ net1076 VGND VPWR _0134_ mac2.products_ff\[74\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5312_ VGND VPWR _2094_ _2096_ _2097_ _2095_ sg13g2_a21oi_1
X_3573_ _0400_ VPWR _0433_ VGND _0397_ _0401_ sg13g2_o21ai_1
X_6292_ net1045 VGND VPWR net334 mac1.sum_lvl3_ff\[1\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_5243_ _2026_ _2006_ _2025_ _2035_ VPWR VGND sg13g2_a21o_1
Xhold19 mac2.sum_lvl1_ff\[47\] VPWR VGND net59 sg13g2_dlygate4sd3_1
X_5174_ _1969_ _1941_ _1967_ VPWR VGND sg13g2_xnor2_1
X_4125_ _0964_ _0959_ _0962_ VPWR VGND sg13g2_xnor2_1
X_4056_ _0865_ _0896_ _0863_ _0898_ VPWR VGND sg13g2_nand3_1
X_3007_ _2604_ net956 net896 VPWR VGND sg13g2_nand2_1
XFILLER_25_857 VPWR VGND sg13g2_decap_4
XFILLER_36_183 VPWR VGND sg13g2_fill_1
X_4958_ _1758_ net854 net785 VPWR VGND sg13g2_nand2_1
X_4889_ _1696_ DP_4.matrix\[6\] net1002 VPWR VGND sg13g2_nand2_1
X_3909_ _0754_ net977 net1004 VPWR VGND sg13g2_nand2_1
XFILLER_0_934 VPWR VGND sg13g2_decap_8
Xfanout1006 net1007 net1006 VPWR VGND sg13g2_buf_8
Xfanout1017 net1021 net1017 VPWR VGND sg13g2_buf_8
Xfanout1028 net1030 net1028 VPWR VGND sg13g2_buf_8
XFILLER_48_905 VPWR VGND sg13g2_decap_8
Xfanout1039 net1040 net1039 VPWR VGND sg13g2_buf_8
XFILLER_28_640 VPWR VGND sg13g2_fill_2
XFILLER_37_1007 VPWR VGND sg13g2_decap_8
XFILLER_42_164 VPWR VGND sg13g2_decap_4
XFILLER_7_577 VPWR VGND sg13g2_fill_1
XFILLER_39_916 VPWR VGND sg13g2_decap_8
XFILLER_47_960 VPWR VGND sg13g2_decap_8
X_5930_ net959 _0188_ VPWR VGND sg13g2_buf_1
X_5861_ net927 net755 _2553_ VPWR VGND sg13g2_nor2_1
XFILLER_34_665 VPWR VGND sg13g2_fill_1
X_4812_ _1621_ _1618_ _1622_ VPWR VGND sg13g2_xor2_1
X_5792_ net809 net825 net779 _2498_ VPWR VGND sg13g2_mux2_1
X_4743_ _1553_ _1554_ _1555_ VPWR VGND sg13g2_nor2_1
XFILLER_30_871 VPWR VGND sg13g2_decap_8
X_6413_ net1089 VGND VPWR net191 mac2.sum_lvl1_ff\[46\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_4674_ _1459_ VPWR _1487_ VGND _1457_ _1460_ sg13g2_o21ai_1
X_3625_ _0456_ VPWR _0484_ VGND _0450_ _0457_ sg13g2_o21ai_1
X_3556_ _0414_ _0415_ _0396_ _0417_ VPWR VGND sg13g2_nand3_1
X_6344_ net1072 VGND VPWR _0138_ mac2.products_ff\[5\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6275_ net1041 VGND VPWR net181 mac1.sum_lvl3_ff\[20\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_5226_ _2019_ _2012_ _2018_ VPWR VGND sg13g2_xnor2_1
X_3487_ _0349_ net992 net925 VPWR VGND sg13g2_nand2_1
XFILLER_29_426 VPWR VGND sg13g2_fill_1
X_5157_ _1951_ _1943_ _1952_ VPWR VGND sg13g2_nor2b_1
X_4108_ _0948_ _0933_ _0947_ VPWR VGND sg13g2_nand2_1
X_5088_ _1873_ VPWR _1885_ VGND _1881_ _1883_ sg13g2_o21ai_1
X_4039_ _0881_ _0875_ _0880_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_337 VPWR VGND sg13g2_fill_1
XFILLER_21_860 VPWR VGND sg13g2_fill_1
XFILLER_43_1011 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_757 VPWR VGND sg13g2_decap_8
XFILLER_29_993 VPWR VGND sg13g2_decap_8
XFILLER_16_643 VPWR VGND sg13g2_fill_2
XFILLER_44_963 VPWR VGND sg13g2_decap_8
XFILLER_16_654 VPWR VGND sg13g2_fill_1
XFILLER_43_495 VPWR VGND sg13g2_fill_1
XFILLER_31_624 VPWR VGND sg13g2_fill_2
XFILLER_12_860 VPWR VGND sg13g2_fill_2
Xhold308 _2301_ VPWR VGND net348 sg13g2_dlygate4sd3_1
X_3410_ net935 net987 net939 _0275_ VPWR VGND net985 sg13g2_nand4_1
Xhold319 DP_4.matrix\[1\] VPWR VGND net359 sg13g2_dlygate4sd3_1
X_4390_ _1189_ VPWR _1217_ VGND _1183_ _1190_ sg13g2_o21ai_1
X_3341_ _2928_ _2913_ _2927_ VPWR VGND sg13g2_nand2_1
X_6060_ net1046 VGND VPWR _0193_ DP_1.matrix\[77\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_3272_ _2861_ _2855_ _2860_ VPWR VGND sg13g2_xnor2_1
X_5011_ _1807_ _1806_ _1789_ _1810_ VPWR VGND sg13g2_a21o_1
XFILLER_39_757 VPWR VGND sg13g2_fill_1
XFILLER_38_256 VPWR VGND sg13g2_fill_1
X_5913_ _2585_ VPWR _0251_ VGND _2527_ _2586_ sg13g2_o21ai_1
XFILLER_34_440 VPWR VGND sg13g2_fill_1
XFILLER_35_985 VPWR VGND sg13g2_decap_8
X_5844_ _2542_ net979 net756 VPWR VGND sg13g2_nand2b_1
XFILLER_21_145 VPWR VGND sg13g2_fill_1
X_2987_ VPWR DP_3.I_range.data_plus_4\[6\] net16 VGND sg13g2_inv_1
X_5775_ _2479_ VPWR _2482_ VGND _2480_ _2481_ sg13g2_o21ai_1
X_4726_ VGND VPWR _1538_ _1536_ _1490_ sg13g2_or2_1
X_4657_ VGND VPWR _1467_ _1468_ _1471_ _1462_ sg13g2_a21oi_1
X_3608_ _0468_ _0421_ _0424_ _0465_ VPWR VGND sg13g2_and3_1
X_6327_ net1012 VGND VPWR net355 mac1.total_sum\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4588_ _1401_ _1402_ _1396_ _1404_ VPWR VGND sg13g2_nand3_1
X_3539_ VGND VPWR _0400_ _0398_ _0357_ sg13g2_or2_1
X_6258_ net1047 VGND VPWR net102 mac1.sum_lvl1_ff\[87\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_6189_ net1080 VGND VPWR net135 mac1.sum_lvl2_ff\[10\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5209_ _1968_ _2001_ _1966_ _2003_ VPWR VGND sg13g2_nand3_1
XFILLER_29_245 VPWR VGND sg13g2_fill_2
XFILLER_26_985 VPWR VGND sg13g2_decap_8
XFILLER_41_955 VPWR VGND sg13g2_decap_8
XFILLER_5_812 VPWR VGND sg13g2_decap_8
XFILLER_5_878 VPWR VGND sg13g2_fill_2
XFILLER_36_705 VPWR VGND sg13g2_fill_1
XFILLER_17_996 VPWR VGND sg13g2_decap_8
X_3890_ _0733_ _0734_ _0728_ _0736_ VPWR VGND sg13g2_nand3_1
XFILLER_32_955 VPWR VGND sg13g2_decap_8
X_5560_ _2285_ _2280_ _2284_ _2290_ VPWR VGND sg13g2_a21o_1
X_4511_ _1332_ _1331_ _1334_ VPWR VGND sg13g2_xor2_1
X_5491_ _2237_ net511 mac2.sum_lvl2_ff\[12\] VPWR VGND sg13g2_nand2_1
Xhold116 mac2.sum_lvl1_ff\[43\] VPWR VGND net156 sg13g2_dlygate4sd3_1
Xhold105 mac2.sum_lvl2_ff\[39\] VPWR VGND net145 sg13g2_dlygate4sd3_1
X_4442_ VGND VPWR _1236_ _1239_ _1268_ _1234_ sg13g2_a21oi_1
Xhold138 mac2.sum_lvl1_ff\[14\] VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold149 mac2.products_ff\[75\] VPWR VGND net189 sg13g2_dlygate4sd3_1
Xhold127 mac2.products_ff\[80\] VPWR VGND net167 sg13g2_dlygate4sd3_1
X_4373_ _1201_ _1155_ _1158_ _1198_ VPWR VGND sg13g2_and3_1
X_6112_ net1067 VGND VPWR net64 mac1.sum_lvl1_ff\[5\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3324_ _2910_ _2906_ _0097_ VPWR VGND sg13g2_xor2_1
X_6043_ net1079 VGND VPWR _0180_ DP_1.matrix\[36\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_3255_ _2845_ _2817_ _2844_ VPWR VGND sg13g2_nand2_1
X_3186_ _2740_ VPWR _2777_ VGND _2698_ _2741_ sg13g2_o21ai_1
X_5827_ VGND VPWR net754 _2530_ _0173_ _2529_ sg13g2_a21oi_1
XFILLER_23_977 VPWR VGND sg13g2_decap_8
XFILLER_22_487 VPWR VGND sg13g2_fill_2
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
X_5758_ VGND VPWR net869 net767 _2465_ net780 sg13g2_a21oi_1
X_4709_ _1520_ _1521_ _1486_ _1522_ VPWR VGND sg13g2_nand3_1
X_5689_ net772 VPWR _2398_ VGND net970 net773 sg13g2_o21ai_1
XFILLER_40_1025 VPWR VGND sg13g2_decap_4
XFILLER_43_73 VPWR VGND sg13g2_decap_4
XFILLER_9_403 VPWR VGND sg13g2_fill_1
XFILLER_14_999 VPWR VGND sg13g2_decap_8
XFILLER_13_498 VPWR VGND sg13g2_decap_4
XFILLER_4_78 VPWR VGND sg13g2_fill_1
XFILLER_1_892 VPWR VGND sg13g2_decap_8
XFILLER_49_863 VPWR VGND sg13g2_decap_8
X_3040_ _2627_ VPWR _2635_ VGND _2619_ _2629_ sg13g2_o21ai_1
XFILLER_36_502 VPWR VGND sg13g2_fill_1
XFILLER_36_524 VPWR VGND sg13g2_decap_4
XFILLER_36_535 VPWR VGND sg13g2_decap_4
X_4991_ _1790_ net852 net785 VPWR VGND sg13g2_nand2_1
X_3942_ _0762_ VPWR _0787_ VGND _0783_ _0785_ sg13g2_o21ai_1
X_3873_ _0716_ _0718_ _0719_ VPWR VGND sg13g2_nor2b_1
X_5612_ VGND VPWR _2325_ _2327_ _2330_ _2329_ sg13g2_a21oi_1
X_5543_ _2275_ net438 _0062_ VPWR VGND sg13g2_nor2b_1
X_5474_ mac2.sum_lvl2_ff\[28\] mac2.sum_lvl2_ff\[9\] _2223_ VPWR VGND sg13g2_nor2_1
X_4425_ _1251_ net866 net995 VPWR VGND sg13g2_nand2_1
X_4356_ _1141_ VPWR _1184_ VGND _1139_ _1142_ sg13g2_o21ai_1
X_3307_ _2895_ _2888_ _2894_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_1009 VPWR VGND sg13g2_decap_8
X_4287_ _1078_ VPWR _1117_ VGND _1079_ _1080_ sg13g2_o21ai_1
X_3238_ _2827_ _2819_ _2828_ VPWR VGND sg13g2_nor2b_1
X_6026_ net1065 VGND VPWR _0163_ DP_2.matrix\[8\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3169_ _2750_ _2758_ _2760_ _2761_ VPWR VGND sg13g2_or3_1
XFILLER_7_929 VPWR VGND sg13g2_decap_8
Xhold480 _2162_ VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold491 mac2.sum_lvl2_ff\[15\] VPWR VGND net531 sg13g2_dlygate4sd3_1
Xfanout960 net961 net960 VPWR VGND sg13g2_buf_2
Xfanout993 net358 net993 VPWR VGND sg13g2_buf_8
Xfanout971 net972 net971 VPWR VGND sg13g2_buf_8
Xfanout982 net502 net982 VPWR VGND sg13g2_buf_8
XFILLER_38_62 VPWR VGND sg13g2_fill_2
XFILLER_6_940 VPWR VGND sg13g2_decap_8
Xclkload14 VPWR clkload14/Y clknet_leaf_66_clk VGND sg13g2_inv_1
XFILLER_47_1009 VPWR VGND sg13g2_decap_8
X_4210_ _1040_ _1039_ _1022_ _1042_ VPWR VGND sg13g2_a21o_1
X_5190_ _1984_ _1978_ _1983_ VPWR VGND sg13g2_xnor2_1
X_4141_ _0979_ _0966_ _0978_ VPWR VGND sg13g2_xnor2_1
X_4072_ _0910_ _0912_ _0913_ VPWR VGND sg13g2_nor2_1
X_3023_ VGND VPWR _2619_ _2618_ _2616_ sg13g2_or2_1
XFILLER_37_844 VPWR VGND sg13g2_fill_2
XFILLER_36_332 VPWR VGND sg13g2_fill_2
XFILLER_37_888 VPWR VGND sg13g2_decap_8
XFILLER_24_538 VPWR VGND sg13g2_fill_1
X_4974_ _1763_ _1771_ _1773_ _1774_ VPWR VGND sg13g2_or3_1
X_3925_ _0770_ _0769_ _0768_ VPWR VGND sg13g2_nand2b_1
X_3856_ _0700_ _0699_ _0694_ _0703_ VPWR VGND sg13g2_a21o_1
Xclkload8 clknet_4_11_0_clk clkload8/X VPWR VGND sg13g2_buf_8
X_3787_ _0636_ DP_2.matrix\[40\] net977 net915 net975 VPWR VGND sg13g2_a22oi_1
X_5526_ mac2.sum_lvl3_ff\[25\] net418 _2263_ VPWR VGND sg13g2_nor2_1
X_5457_ _0043_ _2207_ net449 VPWR VGND sg13g2_xnor2_1
X_4408_ _1197_ _1233_ _1195_ _1235_ VPWR VGND sg13g2_nand3_1
X_5388_ _2156_ mac1.sum_lvl3_ff\[26\] net483 VPWR VGND sg13g2_xnor2_1
X_4339_ VGND VPWR _1167_ _1135_ _1133_ sg13g2_or2_1
XFILLER_46_129 VPWR VGND sg13g2_fill_1
X_6009_ net1064 VGND VPWR _0076_ mac1.products_ff\[70\] clknet_leaf_55_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_66_clk clknet_4_0_0_clk clknet_leaf_66_clk VPWR VGND sg13g2_buf_8
XFILLER_27_332 VPWR VGND sg13g2_fill_2
XFILLER_15_516 VPWR VGND sg13g2_fill_2
XFILLER_28_888 VPWR VGND sg13g2_decap_8
XFILLER_3_921 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_fill_1
XFILLER_3_998 VPWR VGND sg13g2_decap_8
XFILLER_49_83 VPWR VGND sg13g2_decap_8
XFILLER_38_608 VPWR VGND sg13g2_fill_2
Xfanout790 net300 net790 VPWR VGND sg13g2_buf_8
XFILLER_46_630 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_57_clk clknet_4_9_0_clk clknet_leaf_57_clk VPWR VGND sg13g2_buf_8
XFILLER_18_332 VPWR VGND sg13g2_fill_1
XFILLER_46_674 VPWR VGND sg13g2_fill_2
XFILLER_34_814 VPWR VGND sg13g2_fill_2
X_3710_ _0548_ _0542_ _0550_ _0566_ VPWR VGND sg13g2_a21o_1
X_4690_ _1498_ VPWR _1503_ VGND _1500_ _1501_ sg13g2_o21ai_1
X_3641_ VGND VPWR _0462_ _0464_ _0500_ _0499_ sg13g2_a21oi_1
X_3572_ _0391_ VPWR _0432_ VGND _0349_ _0389_ sg13g2_o21ai_1
X_6360_ net1073 VGND VPWR _0127_ mac2.products_ff\[73\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5311_ net534 _2094_ _0010_ VPWR VGND sg13g2_xor2_1
X_6291_ net1043 VGND VPWR net266 mac1.sum_lvl3_ff\[0\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_5242_ _2034_ _2030_ _0152_ VPWR VGND sg13g2_xor2_1
X_5173_ _1968_ _1941_ _1967_ VPWR VGND sg13g2_nand2_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
X_4124_ _0963_ _0962_ _0959_ VPWR VGND sg13g2_nand2b_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ VGND VPWR _0863_ _0865_ _0897_ _0896_ sg13g2_a21oi_1
Xclkbuf_leaf_48_clk clknet_4_11_0_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
X_3006_ VGND VPWR _2596_ _2599_ _2603_ _2597_ sg13g2_a21oi_1
XFILLER_25_836 VPWR VGND sg13g2_decap_4
X_4957_ _1749_ VPWR _1757_ VGND _1741_ _1751_ sg13g2_o21ai_1
X_4888_ _1695_ DP_4.matrix\[7\] net1002 VPWR VGND sg13g2_nand2_1
X_3908_ _0725_ VPWR _0753_ VGND _0723_ _0726_ sg13g2_o21ai_1
X_3839_ _0684_ _0683_ _0686_ VPWR VGND sg13g2_xor2_1
XFILLER_20_574 VPWR VGND sg13g2_fill_2
X_6489_ net1026 VGND VPWR net6 DP_1.Q_range.out_data\[3\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5509_ _2250_ mac2.sum_lvl3_ff\[21\] mac2.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_0_913 VPWR VGND sg13g2_decap_8
Xfanout1007 DP_1.matrix\[80\] net1007 VPWR VGND sg13g2_buf_1
Xfanout1018 net1021 net1018 VPWR VGND sg13g2_buf_8
Xfanout1029 net1030 net1029 VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_39_clk clknet_4_14_0_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_27_151 VPWR VGND sg13g2_fill_2
XFILLER_28_674 VPWR VGND sg13g2_decap_8
XFILLER_15_313 VPWR VGND sg13g2_fill_2
XFILLER_16_847 VPWR VGND sg13g2_fill_1
XFILLER_15_346 VPWR VGND sg13g2_fill_2
XFILLER_42_187 VPWR VGND sg13g2_fill_1
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
XFILLER_18_140 VPWR VGND sg13g2_fill_2
X_5860_ VGND VPWR net757 _2552_ _0200_ net432 sg13g2_a21oi_1
XFILLER_34_633 VPWR VGND sg13g2_decap_4
X_4811_ _1621_ _1576_ _1619_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_121 VPWR VGND sg13g2_fill_2
X_5791_ _2494_ VPWR _2497_ VGND _2495_ _2496_ sg13g2_o21ai_1
XFILLER_22_828 VPWR VGND sg13g2_fill_2
X_4742_ _1554_ net1001 net831 net872 net828 VPWR VGND sg13g2_a22oi_1
XFILLER_21_349 VPWR VGND sg13g2_fill_1
X_4673_ _1475_ VPWR _1486_ VGND _1455_ _1476_ sg13g2_o21ai_1
X_3624_ _0481_ _0473_ _0483_ VPWR VGND sg13g2_xor2_1
X_6412_ net1089 VGND VPWR net62 mac2.sum_lvl1_ff\[45\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3555_ _0416_ _0396_ _0414_ _0415_ VPWR VGND sg13g2_and3_1
X_6343_ net1072 VGND VPWR _0088_ mac2.products_ff\[4\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_6274_ net1031 VGND VPWR net199 mac2.sum_lvl1_ff\[87\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3486_ _0348_ net925 net993 net926 net992 VPWR VGND sg13g2_a22oi_1
X_5225_ _2018_ _2013_ _2016_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_5156_ _1951_ _1944_ _1950_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_909 VPWR VGND sg13g2_decap_8
X_4107_ _0947_ _0918_ _0945_ VPWR VGND sg13g2_xnor2_1
X_5087_ _1873_ _1881_ _1883_ _1884_ VPWR VGND sg13g2_or3_1
X_4038_ _0879_ _0876_ _0880_ VPWR VGND sg13g2_xor2_1
XFILLER_24_165 VPWR VGND sg13g2_fill_2
X_5989_ net1033 VGND VPWR DP_3.Q_range.data_plus_4\[6\] DP_3.Q_range.out_data\[5\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_21_850 VPWR VGND sg13g2_fill_2
XFILLER_40_658 VPWR VGND sg13g2_fill_2
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_29_972 VPWR VGND sg13g2_decap_8
XFILLER_35_408 VPWR VGND sg13g2_fill_2
XFILLER_44_942 VPWR VGND sg13g2_decap_8
XFILLER_43_463 VPWR VGND sg13g2_fill_2
XFILLER_12_872 VPWR VGND sg13g2_fill_2
Xhold309 _0053_ VPWR VGND net349 sg13g2_dlygate4sd3_1
X_3340_ _2927_ _2898_ _2925_ VPWR VGND sg13g2_xnor2_1
X_3271_ _2859_ _2856_ _2860_ VPWR VGND sg13g2_xor2_1
X_5010_ VGND VPWR _1806_ _1807_ _1809_ _1789_ sg13g2_a21oi_1
XFILLER_38_202 VPWR VGND sg13g2_fill_1
X_5912_ _2521_ _2523_ _2586_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_964 VPWR VGND sg13g2_decap_8
X_5843_ VGND VPWR net756 _2541_ _0178_ _2540_ sg13g2_a21oi_1
XFILLER_10_809 VPWR VGND sg13g2_fill_2
XFILLER_22_658 VPWR VGND sg13g2_fill_1
X_5774_ net769 VPWR _2481_ VGND net874 net777 sg13g2_o21ai_1
X_2986_ VPWR DP_1.I_range.data_plus_4\[6\] net4 VGND sg13g2_inv_1
X_4725_ _1537_ net881 net821 VPWR VGND sg13g2_nand2_1
X_4656_ _1467_ _1468_ _1462_ _1470_ VPWR VGND sg13g2_nand3_1
X_3607_ _0424_ _0421_ _0465_ _0467_ VPWR VGND sg13g2_a21o_1
X_4587_ _1403_ _1396_ _1401_ _1402_ VPWR VGND sg13g2_and3_1
X_6326_ net1012 VGND VPWR net385 mac1.total_sum\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3538_ _0399_ net929 net984 VPWR VGND sg13g2_nand2_1
X_3469_ _0327_ VPWR _0332_ VGND _0328_ _0330_ sg13g2_o21ai_1
X_6257_ net1042 VGND VPWR net206 mac1.sum_lvl1_ff\[86\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6188_ net1080 VGND VPWR net71 mac1.sum_lvl2_ff\[9\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5208_ VGND VPWR _1966_ _1968_ _2002_ _2001_ sg13g2_a21oi_1
XFILLER_18_909 VPWR VGND sg13g2_fill_1
X_5139_ _1933_ _1900_ _1935_ VPWR VGND sg13g2_xor2_1
XFILLER_45_706 VPWR VGND sg13g2_fill_2
XFILLER_45_739 VPWR VGND sg13g2_fill_1
XFILLER_44_216 VPWR VGND sg13g2_fill_2
XFILLER_26_964 VPWR VGND sg13g2_decap_8
XFILLER_13_625 VPWR VGND sg13g2_fill_2
XFILLER_41_934 VPWR VGND sg13g2_decap_8
XFILLER_13_636 VPWR VGND sg13g2_fill_1
XFILLER_13_658 VPWR VGND sg13g2_decap_8
XFILLER_9_629 VPWR VGND sg13g2_fill_2
XFILLER_12_157 VPWR VGND sg13g2_decap_4
XFILLER_13_669 VPWR VGND sg13g2_fill_1
XFILLER_48_500 VPWR VGND sg13g2_fill_2
XFILLER_35_205 VPWR VGND sg13g2_fill_1
XFILLER_35_216 VPWR VGND sg13g2_fill_1
XFILLER_17_975 VPWR VGND sg13g2_decap_8
XFILLER_32_934 VPWR VGND sg13g2_decap_8
XFILLER_12_691 VPWR VGND sg13g2_fill_2
X_4510_ _1333_ _1331_ _1332_ VPWR VGND sg13g2_nand2_1
XFILLER_11_190 VPWR VGND sg13g2_fill_1
X_5490_ _2234_ _2235_ _2236_ VPWR VGND sg13g2_nor2_1
XFILLER_7_161 VPWR VGND sg13g2_fill_1
Xhold106 mac1.sum_lvl1_ff\[0\] VPWR VGND net146 sg13g2_dlygate4sd3_1
Xhold117 mac1.sum_lvl1_ff\[5\] VPWR VGND net157 sg13g2_dlygate4sd3_1
X_4441_ _1265_ _1266_ _1267_ VPWR VGND sg13g2_nor2b_1
Xhold128 mac2.products_ff\[83\] VPWR VGND net168 sg13g2_dlygate4sd3_1
Xhold139 mac1.products_ff\[13\] VPWR VGND net179 sg13g2_dlygate4sd3_1
X_6111_ net1075 VGND VPWR _0227_ DP_3.matrix\[7\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_4372_ _1158_ _1155_ _1198_ _1200_ VPWR VGND sg13g2_a21o_1
X_3323_ _2911_ _2906_ _2910_ VPWR VGND sg13g2_nand2_1
X_3254_ _2842_ _2818_ _2844_ VPWR VGND sg13g2_xor2_1
X_6042_ net1065 VGND VPWR _0179_ DP_1.matrix\[7\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_39_500 VPWR VGND sg13g2_decap_4
XFILLER_39_533 VPWR VGND sg13g2_decap_8
X_3185_ _0103_ _2731_ _2775_ VPWR VGND sg13g2_xnor2_1
XFILLER_42_709 VPWR VGND sg13g2_fill_2
XFILLER_26_249 VPWR VGND sg13g2_fill_1
X_5826_ _2388_ _2384_ _2530_ VPWR VGND sg13g2_xor2_1
XFILLER_33_1000 VPWR VGND sg13g2_decap_8
X_5757_ net884 _2463_ _2464_ VPWR VGND sg13g2_nor2_1
X_4708_ _1496_ VPWR _1521_ VGND _1517_ _1519_ sg13g2_o21ai_1
X_5688_ net985 net775 _2397_ VPWR VGND sg13g2_nor2_1
X_4639_ _1450_ _1452_ _1453_ VPWR VGND sg13g2_nor2b_1
X_6309_ net1058 VGND VPWR net169 mac2.sum_lvl3_ff\[22\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_40_1004 VPWR VGND sg13g2_decap_8
XFILLER_45_558 VPWR VGND sg13g2_fill_1
XFILLER_14_978 VPWR VGND sg13g2_decap_8
XFILLER_43_85 VPWR VGND sg13g2_fill_1
X_4990_ _1772_ VPWR _1789_ VGND _1763_ _1773_ sg13g2_o21ai_1
XFILLER_44_591 VPWR VGND sg13g2_decap_4
X_3941_ _0762_ _0783_ _0785_ _0786_ VPWR VGND sg13g2_or3_1
XFILLER_17_794 VPWR VGND sg13g2_fill_1
X_3872_ VGND VPWR _0718_ _0717_ _0684_ sg13g2_or2_1
XFILLER_17_1017 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
X_5611_ _2329_ mac1.total_sum\[8\] mac2.total_sum\[8\] VPWR VGND sg13g2_xnor2_1
X_5542_ _2272_ _2274_ net437 _2276_ VPWR VGND sg13g2_nand3_1
XFILLER_8_470 VPWR VGND sg13g2_fill_1
X_5473_ VGND VPWR mac2.sum_lvl2_ff\[27\] mac2.sum_lvl2_ff\[8\] _2222_ _2220_ sg13g2_a21oi_1
X_4424_ VGND VPWR _1250_ _1223_ _1221_ sg13g2_or2_1
X_4355_ _1183_ _1178_ _1182_ VPWR VGND sg13g2_xnor2_1
X_3306_ _2894_ _2889_ _2892_ VPWR VGND sg13g2_xnor2_1
X_4286_ _1115_ _1052_ _1116_ VPWR VGND sg13g2_xor2_1
X_3237_ _2827_ _2820_ _2826_ VPWR VGND sg13g2_xnor2_1
X_6025_ net1046 VGND VPWR _0162_ DP_1.matrix\[80\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_3168_ VGND VPWR _2756_ _2757_ _2760_ _2751_ sg13g2_a21oi_1
XFILLER_42_506 VPWR VGND sg13g2_fill_2
X_3099_ VGND VPWR _2634_ _2660_ _2693_ _2659_ sg13g2_a21oi_1
X_5809_ _2515_ _2514_ _2510_ VPWR VGND sg13g2_nand2b_1
Xhold481 _0029_ VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold470 DP_1.matrix\[4\] VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold492 _2248_ VPWR VGND net532 sg13g2_dlygate4sd3_1
Xfanout950 net951 net950 VPWR VGND sg13g2_buf_1
Xfanout961 net962 net961 VPWR VGND sg13g2_buf_8
Xfanout994 DP_4.matrix\[80\] net994 VPWR VGND sg13g2_buf_8
Xfanout972 net491 net972 VPWR VGND sg13g2_buf_8
Xfanout983 net984 net983 VPWR VGND sg13g2_buf_8
XFILLER_46_812 VPWR VGND sg13g2_fill_2
XFILLER_18_536 VPWR VGND sg13g2_fill_1
XFILLER_46_889 VPWR VGND sg13g2_decap_8
XFILLER_41_550 VPWR VGND sg13g2_decap_8
XFILLER_41_561 VPWR VGND sg13g2_fill_2
Xclkload15 VPWR clkload15/Y clknet_leaf_28_clk VGND sg13g2_inv_1
XFILLER_10_992 VPWR VGND sg13g2_decap_8
XFILLER_6_996 VPWR VGND sg13g2_decap_8
X_4140_ _0978_ _0975_ _0977_ VPWR VGND sg13g2_xnor2_1
X_4071_ _0912_ net906 net966 net908 net964 VPWR VGND sg13g2_a22oi_1
XFILLER_48_160 VPWR VGND sg13g2_fill_2
X_3022_ _2602_ _2617_ _2618_ VPWR VGND sg13g2_nor2_1
XFILLER_37_867 VPWR VGND sg13g2_decap_8
X_4973_ VGND VPWR _1769_ _1770_ _1773_ _1764_ sg13g2_a21oi_1
X_3924_ _0764_ VPWR _0769_ VGND _0766_ _0767_ sg13g2_o21ai_1
X_3855_ _0699_ _0700_ _0694_ _0702_ VPWR VGND sg13g2_nand3_1
Xclkload9 clknet_4_12_0_clk clkload9/X VPWR VGND sg13g2_buf_8
X_3786_ _0077_ _0621_ _0634_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_1025 VPWR VGND sg13g2_decap_4
X_5525_ VGND VPWR _2259_ _2261_ _2262_ _2260_ sg13g2_a21oi_1
X_5456_ net448 mac2.sum_lvl2_ff\[24\] _2209_ VPWR VGND sg13g2_xor2_1
X_4407_ VGND VPWR _1195_ _1197_ _1234_ _1233_ sg13g2_a21oi_1
X_5387_ mac1.sum_lvl3_ff\[26\] net483 _2155_ VPWR VGND sg13g2_and2_1
XFILLER_8_1015 VPWR VGND sg13g2_decap_8
X_4338_ _1125_ VPWR _1166_ VGND _1084_ _1123_ sg13g2_o21ai_1
X_4269_ _1099_ net855 DP_4.matrix\[36\] net858 net815 VPWR VGND sg13g2_a22oi_1
X_6008_ net1043 VGND VPWR _0075_ mac1.products_ff\[69\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_28_867 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_fill_1
XFILLER_40_31 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_fill_2
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_8
Xfanout780 _2448_ net780 VPWR VGND sg13g2_buf_8
XFILLER_19_845 VPWR VGND sg13g2_fill_1
XFILLER_46_664 VPWR VGND sg13g2_fill_1
X_3640_ _0499_ _0471_ _0497_ VPWR VGND sg13g2_xnor2_1
X_3571_ _0417_ VPWR _0431_ VGND _0395_ _0418_ sg13g2_o21ai_1
X_5310_ net533 mac1.sum_lvl2_ff\[23\] _2096_ VPWR VGND sg13g2_xor2_1
X_6290_ net1065 VGND VPWR net129 mac1.sum_lvl3_ff\[35\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_5241_ VGND VPWR _2033_ _2034_ _2032_ _1973_ sg13g2_a21oi_2
X_5172_ _1965_ _1942_ _1967_ VPWR VGND sg13g2_xor2_1
X_4123_ _0961_ _0936_ _0962_ VPWR VGND sg13g2_xor2_1
X_4054_ _0894_ _0873_ _0896_ VPWR VGND sg13g2_xor2_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
X_3005_ _2602_ net958 net894 VPWR VGND sg13g2_nand2_1
XFILLER_24_336 VPWR VGND sg13g2_fill_1
X_4956_ _1755_ _1737_ _0093_ VPWR VGND sg13g2_xor2_1
XFILLER_33_881 VPWR VGND sg13g2_decap_8
X_4887_ _1694_ net875 DP_4.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_3907_ _0741_ VPWR _0752_ VGND _0721_ _0742_ sg13g2_o21ai_1
X_3838_ _0685_ _0683_ _0684_ VPWR VGND sg13g2_nand2b_1
XFILLER_3_218 VPWR VGND sg13g2_fill_1
X_3769_ _0619_ _0616_ _0620_ VPWR VGND sg13g2_xor2_1
X_5508_ _2249_ net474 net305 VPWR VGND sg13g2_nand2_1
X_6488_ net1027 VGND VPWR net5 DP_1.Q_range.out_data\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5439_ mac2.sum_lvl2_ff\[20\] mac2.sum_lvl2_ff\[1\] _2196_ VPWR VGND sg13g2_nor2_1
Xfanout1019 net1020 net1019 VPWR VGND sg13g2_buf_8
Xfanout1008 net1009 net1008 VPWR VGND sg13g2_buf_8
XFILLER_0_969 VPWR VGND sg13g2_decap_8
XFILLER_27_141 VPWR VGND sg13g2_fill_1
XFILLER_11_564 VPWR VGND sg13g2_fill_2
XFILLER_47_995 VPWR VGND sg13g2_decap_8
X_4810_ VGND VPWR _1620_ _1619_ _1576_ sg13g2_or2_1
X_5790_ net768 VPWR _2496_ VGND net822 net777 sg13g2_o21ai_1
XFILLER_15_881 VPWR VGND sg13g2_fill_1
X_4741_ net832 net828 net872 net1002 _1553_ VPWR VGND sg13g2_and4_1
XFILLER_21_339 VPWR VGND sg13g2_fill_2
X_4672_ _1484_ _1483_ _0146_ VPWR VGND sg13g2_xor2_1
X_3623_ _0481_ _0473_ _0482_ VPWR VGND sg13g2_nor2b_1
X_6411_ net1088 VGND VPWR net186 mac2.sum_lvl1_ff\[44\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3554_ _0403_ VPWR _0415_ VGND _0411_ _0413_ sg13g2_o21ai_1
X_6342_ net1059 VGND VPWR _0087_ mac2.products_ff\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_3485_ _0324_ VPWR _0347_ VGND _0289_ _0322_ sg13g2_o21ai_1
X_6273_ net1032 VGND VPWR net258 mac2.sum_lvl1_ff\[86\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5224_ _2017_ _2016_ _2013_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_5155_ _1949_ _1945_ _1950_ VPWR VGND sg13g2_xor2_1
X_4106_ _0946_ _0945_ _0918_ VPWR VGND sg13g2_nand2b_1
X_5086_ VGND VPWR _1879_ _1880_ _1883_ _1874_ sg13g2_a21oi_1
X_4037_ _0879_ _0853_ _0877_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_984 VPWR VGND sg13g2_decap_8
XFILLER_25_678 VPWR VGND sg13g2_decap_8
X_5988_ net1033 VGND VPWR net11 DP_3.Q_range.out_data\[4\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_4939_ _1724_ _1739_ _1740_ VPWR VGND sg13g2_nor2_1
XFILLER_40_637 VPWR VGND sg13g2_fill_1
XFILLER_20_361 VPWR VGND sg13g2_fill_1
XFILLER_21_55 VPWR VGND sg13g2_fill_2
XFILLER_21_66 VPWR VGND sg13g2_fill_1
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_29_951 VPWR VGND sg13g2_decap_8
XFILLER_46_85 VPWR VGND sg13g2_decap_4
XFILLER_44_921 VPWR VGND sg13g2_decap_8
XFILLER_16_645 VPWR VGND sg13g2_fill_1
XFILLER_44_998 VPWR VGND sg13g2_decap_8
X_3270_ _2859_ _2833_ _2857_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_4 VPWR VGND sg13g2_fill_2
XFILLER_39_726 VPWR VGND sg13g2_fill_2
XFILLER_38_214 VPWR VGND sg13g2_fill_2
XFILLER_38_247 VPWR VGND sg13g2_fill_2
X_5911_ _2585_ net820 net760 VPWR VGND sg13g2_nand2_1
XFILLER_35_943 VPWR VGND sg13g2_decap_8
X_5842_ _2403_ _2401_ _2541_ VPWR VGND sg13g2_xor2_1
X_5773_ net860 net779 _2480_ VPWR VGND sg13g2_nor2_1
X_4724_ _1536_ net881 net820 VPWR VGND sg13g2_nand2_1
X_2985_ VPWR _2589_ DP_3.Q_range.out_data\[5\] VGND sg13g2_inv_1
X_4655_ _1469_ _1462_ _1467_ _1468_ VPWR VGND sg13g2_and3_1
X_3606_ VGND VPWR _0421_ _0424_ _0466_ _0465_ sg13g2_a21oi_1
X_4586_ _1397_ VPWR _1402_ VGND _1398_ _1400_ sg13g2_o21ai_1
X_6325_ net1012 VGND VPWR net435 mac1.total_sum\[2\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3537_ _0398_ net928 net984 VPWR VGND sg13g2_nand2_1
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
X_3468_ _0327_ _0328_ _0330_ _0331_ VPWR VGND sg13g2_or3_1
X_6256_ net1049 VGND VPWR net44 mac1.sum_lvl1_ff\[85\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3399_ _2980_ _2979_ _2969_ VPWR VGND sg13g2_nand2b_1
X_6187_ net1080 VGND VPWR net151 mac1.sum_lvl2_ff\[8\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5207_ _1999_ _1976_ _2001_ VPWR VGND sg13g2_xor2_1
X_5138_ _1934_ _1900_ _1933_ VPWR VGND sg13g2_nand2b_1
XFILLER_45_729 VPWR VGND sg13g2_fill_2
X_5069_ _1839_ VPWR _1866_ VGND _1830_ _1840_ sg13g2_o21ai_1
XFILLER_26_943 VPWR VGND sg13g2_decap_8
XFILLER_25_486 VPWR VGND sg13g2_fill_1
XFILLER_41_913 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_fill_1
XFILLER_17_954 VPWR VGND sg13g2_decap_8
XFILLER_32_913 VPWR VGND sg13g2_decap_8
XFILLER_8_630 VPWR VGND sg13g2_decap_8
XFILLER_40_990 VPWR VGND sg13g2_decap_8
Xhold107 mac1.products_ff\[6\] VPWR VGND net147 sg13g2_dlygate4sd3_1
X_4440_ _1232_ _1264_ _1230_ _1266_ VPWR VGND sg13g2_nand3_1
Xhold118 mac1.sum_lvl2_ff\[51\] VPWR VGND net158 sg13g2_dlygate4sd3_1
Xhold129 mac2.sum_lvl2_ff\[40\] VPWR VGND net169 sg13g2_dlygate4sd3_1
X_6110_ net1075 VGND VPWR _0226_ DP_3.matrix\[6\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_4371_ VGND VPWR _1155_ _1158_ _1199_ _1198_ sg13g2_a21oi_1
X_3322_ VGND VPWR _2909_ _2910_ _2908_ _2850_ sg13g2_a21oi_2
X_3253_ _2843_ _2818_ _2842_ VPWR VGND sg13g2_nand2_1
X_6041_ net1065 VGND VPWR _0178_ DP_1.matrix\[6\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3184_ _2730_ _2775_ _2729_ _2776_ VPWR VGND sg13g2_nand3_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
XFILLER_23_902 VPWR VGND sg13g2_fill_2
X_5825_ net991 net754 _2529_ VPWR VGND sg13g2_nor2_1
XFILLER_22_456 VPWR VGND sg13g2_fill_2
X_5756_ _2463_ _2446_ net780 VPWR VGND sg13g2_nand2_1
XFILLER_31_990 VPWR VGND sg13g2_decap_8
X_5687_ _2396_ net951 net763 VPWR VGND sg13g2_nand2_1
X_4707_ _1496_ _1517_ _1519_ _1520_ VPWR VGND sg13g2_or3_1
X_4638_ VGND VPWR _1452_ _1451_ _1418_ sg13g2_or2_1
XFILLER_2_806 VPWR VGND sg13g2_fill_2
XFILLER_2_817 VPWR VGND sg13g2_decap_4
X_4569_ _1386_ _1384_ _1385_ VPWR VGND sg13g2_nand2_1
X_6308_ net1051 VGND VPWR net145 mac2.sum_lvl3_ff\[21\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_6239_ net1038 VGND VPWR net128 mac2.sum_lvl2_ff\[50\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_13_401 VPWR VGND sg13g2_fill_2
XFILLER_14_902 VPWR VGND sg13g2_decap_4
XFILLER_14_957 VPWR VGND sg13g2_decap_8
XFILLER_25_272 VPWR VGND sg13g2_fill_2
XFILLER_13_445 VPWR VGND sg13g2_fill_2
XFILLER_22_990 VPWR VGND sg13g2_decap_8
XFILLER_49_898 VPWR VGND sg13g2_decap_8
X_3940_ VGND VPWR _0781_ _0782_ _0785_ _0763_ sg13g2_a21oi_1
X_3871_ _0717_ net976 net906 VPWR VGND sg13g2_nand2_1
XFILLER_20_916 VPWR VGND sg13g2_decap_8
X_5610_ _2327_ _2328_ net32 VPWR VGND sg13g2_and2_1
X_5541_ VGND VPWR net437 _2272_ _2275_ _2274_ sg13g2_a21oi_1
XFILLER_9_994 VPWR VGND sg13g2_decap_8
X_5472_ _2220_ _2221_ _0046_ VPWR VGND sg13g2_nor2b_2
X_4423_ _1211_ VPWR _1249_ VGND _1208_ _1212_ sg13g2_o21ai_1
X_4354_ _1182_ _1132_ _1179_ VPWR VGND sg13g2_xnor2_1
X_3305_ _2893_ _2892_ _2889_ VPWR VGND sg13g2_nand2b_1
X_6024_ net1081 VGND VPWR _0161_ DP_1.matrix\[44\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_4285_ _1115_ _1112_ _1114_ VPWR VGND sg13g2_nand2_1
X_3236_ _2825_ _2821_ _2826_ VPWR VGND sg13g2_xor2_1
X_3167_ _2756_ _2757_ _2751_ _2759_ VPWR VGND sg13g2_nand3_1
X_3098_ _2690_ _2662_ _2692_ VPWR VGND sg13g2_xor2_1
X_5808_ _2511_ VPWR _2514_ VGND _2512_ _2513_ sg13g2_o21ai_1
XFILLER_11_949 VPWR VGND sg13g2_decap_8
XFILLER_22_297 VPWR VGND sg13g2_fill_1
X_5739_ DP_3.Q_range.out_data\[3\] DP_3.I_range.out_data\[3\] _2446_ VPWR VGND sg13g2_xor2_1
Xhold460 _2105_ VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold471 mac2.sum_lvl2_ff\[31\] VPWR VGND net511 sg13g2_dlygate4sd3_1
Xhold482 DP_1.matrix\[41\] VPWR VGND net522 sg13g2_dlygate4sd3_1
Xhold493 mac1.sum_lvl2_ff\[4\] VPWR VGND net533 sg13g2_dlygate4sd3_1
XFILLER_49_117 VPWR VGND sg13g2_decap_8
Xfanout951 net297 net951 VPWR VGND sg13g2_buf_8
Xfanout940 net427 net940 VPWR VGND sg13g2_buf_1
Xfanout995 DP_4.matrix\[44\] net995 VPWR VGND sg13g2_buf_8
Xfanout973 DP_1.matrix\[38\] net973 VPWR VGND sg13g2_buf_8
Xfanout984 net503 net984 VPWR VGND sg13g2_buf_8
Xfanout962 net477 net962 VPWR VGND sg13g2_buf_8
XFILLER_46_868 VPWR VGND sg13g2_decap_8
XFILLER_45_334 VPWR VGND sg13g2_fill_1
XFILLER_13_297 VPWR VGND sg13g2_fill_2
XFILLER_9_279 VPWR VGND sg13g2_fill_2
XFILLER_10_971 VPWR VGND sg13g2_decap_8
Xclkload16 VPWR clkload16/Y clknet_leaf_27_clk VGND sg13g2_inv_1
XFILLER_6_975 VPWR VGND sg13g2_decap_8
XFILLER_5_463 VPWR VGND sg13g2_fill_2
X_4070_ VGND VPWR _0911_ _0909_ _0885_ sg13g2_or2_1
X_3021_ _2617_ net956 net892 VPWR VGND sg13g2_nand2_1
XFILLER_37_846 VPWR VGND sg13g2_fill_1
XFILLER_24_529 VPWR VGND sg13g2_decap_8
X_4972_ _1769_ _1770_ _1764_ _1772_ VPWR VGND sg13g2_nand3_1
X_3923_ _0764_ _0766_ _0767_ _0768_ VPWR VGND sg13g2_nor3_1
X_3854_ _0701_ _0694_ _0699_ _0700_ VPWR VGND sg13g2_and3_1
XFILLER_32_584 VPWR VGND sg13g2_fill_2
X_3785_ _0621_ _0634_ _0635_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_1004 VPWR VGND sg13g2_decap_8
X_5524_ net455 _2259_ _0058_ VPWR VGND sg13g2_xor2_1
X_5455_ mac2.sum_lvl2_ff\[24\] net448 _2208_ VPWR VGND sg13g2_nor2_1
X_4406_ _1233_ _1204_ _1231_ VPWR VGND sg13g2_xnor2_1
X_5386_ _0027_ _2152_ net318 VPWR VGND sg13g2_xnor2_1
X_4337_ _1151_ VPWR _1165_ VGND _1129_ _1152_ sg13g2_o21ai_1
X_4268_ net814 net858 net817 _1098_ VPWR VGND net855 sg13g2_nand4_1
X_6007_ net1043 VGND VPWR _0074_ mac1.products_ff\[68\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3219_ _2810_ _2777_ _2809_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_802 VPWR VGND sg13g2_decap_4
XFILLER_39_161 VPWR VGND sg13g2_fill_1
XFILLER_27_334 VPWR VGND sg13g2_fill_1
X_4199_ net818 net816 net863 net862 _1031_ VPWR VGND sg13g2_and4_1
XFILLER_27_356 VPWR VGND sg13g2_fill_2
XFILLER_42_337 VPWR VGND sg13g2_fill_1
XFILLER_3_956 VPWR VGND sg13g2_decap_8
XFILLER_46_1022 VPWR VGND sg13g2_decap_8
Xhold290 DP_4.matrix\[37\] VPWR VGND net330 sg13g2_dlygate4sd3_1
Xfanout792 net303 net792 VPWR VGND sg13g2_buf_8
Xfanout781 net782 net781 VPWR VGND sg13g2_buf_8
Xfanout770 net772 net770 VPWR VGND sg13g2_buf_8
XFILLER_46_676 VPWR VGND sg13g2_fill_1
XFILLER_34_816 VPWR VGND sg13g2_fill_1
XFILLER_42_882 VPWR VGND sg13g2_decap_8
X_3570_ _0393_ VPWR _0430_ VGND _0350_ _0394_ sg13g2_o21ai_1
X_5240_ _2003_ VPWR _2033_ VGND _1971_ _2002_ sg13g2_o21ai_1
X_5171_ _1966_ _1942_ _1965_ VPWR VGND sg13g2_nand2_1
XFILLER_39_2 VPWR VGND sg13g2_fill_1
X_4122_ _0961_ net909 net1008 VPWR VGND sg13g2_nand2_1
X_4053_ _0894_ _0873_ _0895_ VPWR VGND sg13g2_nor2b_1
X_3004_ _2600_ _2594_ _0066_ VPWR VGND sg13g2_xor2_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
X_4955_ _1737_ _1755_ _1756_ VPWR VGND sg13g2_and2_1
X_3906_ _0750_ _0749_ _0124_ VPWR VGND sg13g2_xor2_1
X_4886_ _1677_ _1669_ _1676_ _1693_ VPWR VGND sg13g2_a21o_1
XFILLER_20_532 VPWR VGND sg13g2_fill_2
X_3837_ _0684_ net977 net908 VPWR VGND sg13g2_nand2_1
X_3768_ _0617_ _0618_ _0619_ VPWR VGND sg13g2_nor2_1
XFILLER_3_208 VPWR VGND sg13g2_fill_1
X_5507_ net267 mac2.sum_lvl2_ff\[19\] _0032_ VPWR VGND sg13g2_xor2_1
X_3699_ _0556_ _0553_ _0554_ VPWR VGND sg13g2_xnor2_1
X_6487_ net1020 VGND VPWR net369 mac2.total_sum\[15\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5438_ _2195_ mac2.sum_lvl2_ff\[20\] mac2.sum_lvl2_ff\[1\] VPWR VGND sg13g2_nand2_1
X_5369_ mac1.sum_lvl3_ff\[1\] mac1.sum_lvl3_ff\[21\] _2142_ VPWR VGND sg13g2_xor2_1
XFILLER_0_948 VPWR VGND sg13g2_decap_8
Xfanout1009 net403 net1009 VPWR VGND sg13g2_buf_2
XFILLER_48_919 VPWR VGND sg13g2_decap_8
XFILLER_47_407 VPWR VGND sg13g2_fill_2
XFILLER_19_77 VPWR VGND sg13g2_fill_1
XFILLER_27_153 VPWR VGND sg13g2_fill_1
XFILLER_15_337 VPWR VGND sg13g2_decap_4
XFILLER_15_348 VPWR VGND sg13g2_fill_1
XFILLER_30_318 VPWR VGND sg13g2_fill_1
XFILLER_13_1010 VPWR VGND sg13g2_decap_8
XFILLER_3_764 VPWR VGND sg13g2_fill_2
XFILLER_47_974 VPWR VGND sg13g2_decap_8
XFILLER_46_473 VPWR VGND sg13g2_fill_2
XFILLER_33_123 VPWR VGND sg13g2_fill_1
XFILLER_34_679 VPWR VGND sg13g2_fill_2
X_4740_ _1552_ net828 net1001 VPWR VGND sg13g2_nand2_1
X_4671_ _1485_ _1483_ _1484_ VPWR VGND sg13g2_nand2_1
X_3622_ _0481_ _0474_ _0480_ VPWR VGND sg13g2_xnor2_1
X_6410_ net1081 VGND VPWR net189 mac2.sum_lvl1_ff\[43\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_30_885 VPWR VGND sg13g2_decap_8
X_6341_ net1057 VGND VPWR _0086_ mac2.products_ff\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_3553_ _0403_ _0411_ _0413_ _0414_ VPWR VGND sg13g2_or3_1
X_3484_ _0338_ VPWR _0346_ VGND _0318_ _0339_ sg13g2_o21ai_1
X_6272_ net1033 VGND VPWR net219 mac2.sum_lvl1_ff\[85\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5223_ _2015_ _1989_ _2016_ VPWR VGND sg13g2_xor2_1
X_5154_ _1949_ _1905_ _1947_ VPWR VGND sg13g2_xnor2_1
X_4105_ _0943_ _0903_ _0945_ VPWR VGND sg13g2_xor2_1
X_5085_ _1879_ _1880_ _1874_ _1882_ VPWR VGND sg13g2_nand3_1
X_4036_ VGND VPWR _0878_ _0877_ _0853_ sg13g2_or2_1
XFILLER_38_963 VPWR VGND sg13g2_decap_8
XFILLER_25_646 VPWR VGND sg13g2_decap_4
XFILLER_24_167 VPWR VGND sg13g2_fill_1
X_5987_ net1033 VGND VPWR net10 DP_3.Q_range.out_data\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_4938_ _1739_ net852 net788 VPWR VGND sg13g2_nand2_2
X_4869_ _1677_ _1638_ _1675_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_43_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_930 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
XFILLER_44_977 VPWR VGND sg13g2_decap_8
XFILLER_43_465 VPWR VGND sg13g2_fill_1
XFILLER_7_311 VPWR VGND sg13g2_fill_2
XFILLER_7_36 VPWR VGND sg13g2_fill_1
XFILLER_12_885 VPWR VGND sg13g2_fill_2
XFILLER_39_716 VPWR VGND sg13g2_fill_1
X_5910_ _2584_ VPWR _0250_ VGND net760 _2583_ sg13g2_o21ai_1
XFILLER_35_922 VPWR VGND sg13g2_decap_8
X_5841_ net981 net755 _2540_ VPWR VGND sg13g2_nor2_1
XFILLER_34_465 VPWR VGND sg13g2_fill_1
XFILLER_35_999 VPWR VGND sg13g2_decap_8
X_2984_ VPWR _2588_ DP_3.I_range.out_data\[5\] VGND sg13g2_inv_1
X_5772_ _2479_ net843 net765 VPWR VGND sg13g2_nand2_1
X_4723_ _1535_ net885 net996 VPWR VGND sg13g2_nand2_1
X_4654_ _1463_ VPWR _1468_ VGND _1464_ _1466_ sg13g2_o21ai_1
X_3605_ _0463_ _0430_ _0465_ VPWR VGND sg13g2_xor2_1
X_4585_ _1397_ _1398_ _1400_ _1401_ VPWR VGND sg13g2_or3_1
X_6324_ net1013 VGND VPWR net430 mac1.total_sum\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3536_ _0397_ net988 net927 VPWR VGND sg13g2_nand2_1
X_6255_ net1020 VGND VPWR net202 mac1.sum_lvl1_ff\[84\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3467_ _0330_ net981 net938 net983 net933 VPWR VGND sg13g2_a22oi_1
X_5206_ _1999_ _1976_ _2000_ VPWR VGND sg13g2_nor2b_1
X_6186_ net1079 VGND VPWR net127 mac1.sum_lvl2_ff\[7\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3398_ _2979_ _2970_ _2977_ VPWR VGND sg13g2_xnor2_1
X_5137_ _1933_ _1901_ _1931_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_719 VPWR VGND sg13g2_fill_2
XFILLER_45_708 VPWR VGND sg13g2_fill_1
X_5068_ _1865_ _1820_ _1864_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_218 VPWR VGND sg13g2_fill_1
X_4019_ _0861_ _0849_ _0862_ VPWR VGND sg13g2_xor2_1
XFILLER_26_999 VPWR VGND sg13g2_decap_8
XFILLER_9_609 VPWR VGND sg13g2_fill_2
XFILLER_41_969 VPWR VGND sg13g2_decap_8
XFILLER_10_1013 VPWR VGND sg13g2_decap_8
XFILLER_4_336 VPWR VGND sg13g2_fill_2
XFILLER_48_502 VPWR VGND sg13g2_fill_1
XFILLER_48_524 VPWR VGND sg13g2_fill_2
XFILLER_36_719 VPWR VGND sg13g2_decap_8
XFILLER_16_410 VPWR VGND sg13g2_fill_2
XFILLER_43_240 VPWR VGND sg13g2_fill_1
XFILLER_32_969 VPWR VGND sg13g2_decap_8
Xhold108 mac1.sum_lvl1_ff\[72\] VPWR VGND net148 sg13g2_dlygate4sd3_1
Xhold119 mac2.sum_lvl1_ff\[13\] VPWR VGND net159 sg13g2_dlygate4sd3_1
X_4370_ _1196_ _1164_ _1198_ VPWR VGND sg13g2_xor2_1
X_3321_ _2879_ VPWR _2909_ VGND _2848_ _2878_ sg13g2_o21ai_1
X_6040_ net1047 VGND VPWR _0177_ DP_1.matrix\[5\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3252_ _2841_ _2829_ _2842_ VPWR VGND sg13g2_xor2_1
XFILLER_26_1020 VPWR VGND sg13g2_decap_8
X_3183_ _2773_ _2774_ _2775_ VPWR VGND sg13g2_and2_1
X_5824_ net754 net993 _0172_ VPWR VGND sg13g2_xor2_1
X_5755_ _2462_ _2461_ net767 net765 net854 VPWR VGND sg13g2_a22oi_1
X_5686_ _2395_ _2382_ _2394_ VPWR VGND sg13g2_nand2b_1
X_4706_ VGND VPWR _1515_ _1516_ _1519_ _1497_ sg13g2_a21oi_1
X_4637_ _1451_ net885 net820 VPWR VGND sg13g2_nand2_1
X_4568_ _1385_ _1365_ _1367_ VPWR VGND sg13g2_nand2_1
X_4499_ VGND VPWR _1292_ _1317_ _1322_ _1318_ sg13g2_a21oi_1
X_3519_ _0381_ _0378_ _0380_ VPWR VGND sg13g2_nand2_1
X_6307_ net1051 VGND VPWR net256 mac2.sum_lvl3_ff\[20\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6238_ net1029 VGND VPWR net154 mac2.sum_lvl2_ff\[49\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6169_ net1078 VGND VPWR net237 mac1.sum_lvl1_ff\[42\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_45_516 VPWR VGND sg13g2_fill_1
XFILLER_43_54 VPWR VGND sg13g2_fill_1
XFILLER_43_98 VPWR VGND sg13g2_fill_1
XFILLER_40_276 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_20_clk clknet_4_5_0_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_4_144 VPWR VGND sg13g2_fill_2
XFILLER_49_877 VPWR VGND sg13g2_decap_8
XFILLER_1_1011 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_fill_1
X_3870_ _0716_ net906 DP_1.matrix\[36\] net908 net976 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_11_clk clknet_4_9_0_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_5540_ _2274_ mac2.sum_lvl3_ff\[28\] mac2.sum_lvl3_ff\[8\] VPWR VGND sg13g2_xnor2_1
XFILLER_9_973 VPWR VGND sg13g2_decap_8
X_5471_ _2217_ _2219_ net507 _2221_ VPWR VGND sg13g2_nand3_1
X_4422_ _1248_ _1242_ _1247_ VPWR VGND sg13g2_xnor2_1
X_4353_ _1132_ _1179_ _1181_ VPWR VGND sg13g2_and2_1
X_3304_ _2891_ _2865_ _2892_ VPWR VGND sg13g2_xor2_1
X_4284_ _1111_ _1110_ _1081_ _1114_ VPWR VGND sg13g2_a21o_1
X_3235_ _2825_ _2782_ _2823_ VPWR VGND sg13g2_xnor2_1
X_6023_ net1066 VGND VPWR net446 DP_1.matrix\[8\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3166_ _2758_ _2751_ _2756_ _2757_ VPWR VGND sg13g2_and3_1
XFILLER_39_354 VPWR VGND sg13g2_fill_1
X_3097_ _2691_ _2662_ _2690_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_538 VPWR VGND sg13g2_fill_2
XFILLER_35_582 VPWR VGND sg13g2_fill_1
X_5807_ net768 VPWR _2513_ VGND net824 net777 sg13g2_o21ai_1
X_3999_ _0842_ net968 net906 VPWR VGND sg13g2_nand2_1
X_5738_ _2445_ DP_3.I_range.out_data\[2\] DP_3.Q_range.out_data\[2\] VPWR VGND sg13g2_nand2b_1
X_5669_ _2378_ net771 _2377_ net764 net948 VPWR VGND sg13g2_a22oi_1
Xhold461 _0014_ VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold450 DP_2.matrix\[8\] VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold472 _2237_ VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold494 _2096_ VPWR VGND net534 sg13g2_dlygate4sd3_1
XFILLER_1_136 VPWR VGND sg13g2_fill_1
Xhold483 DP_2.matrix\[40\] VPWR VGND net523 sg13g2_dlygate4sd3_1
Xfanout930 net388 net930 VPWR VGND sg13g2_buf_8
Xfanout941 net942 net941 VPWR VGND sg13g2_buf_8
Xfanout952 net953 net952 VPWR VGND sg13g2_buf_8
XFILLER_1_169 VPWR VGND sg13g2_fill_1
Xfanout974 net371 net974 VPWR VGND sg13g2_buf_2
Xfanout963 net965 net963 VPWR VGND sg13g2_buf_8
Xfanout985 net986 net985 VPWR VGND sg13g2_buf_8
Xfanout996 net476 net996 VPWR VGND sg13g2_buf_8
XFILLER_13_243 VPWR VGND sg13g2_fill_2
XFILLER_13_254 VPWR VGND sg13g2_fill_2
XFILLER_10_950 VPWR VGND sg13g2_decap_8
Xclkload17 clkload17/Y clknet_leaf_56_clk VPWR VGND sg13g2_inv_2
XFILLER_6_954 VPWR VGND sg13g2_decap_8
XFILLER_23_1012 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_4_0_0_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
X_3020_ _2616_ net892 net958 net894 net956 VPWR VGND sg13g2_a22oi_1
X_4971_ _1771_ _1764_ _1769_ _1770_ VPWR VGND sg13g2_and3_1
X_3922_ _0767_ net966 net914 net912 net969 VPWR VGND sg13g2_a22oi_1
XFILLER_17_593 VPWR VGND sg13g2_fill_2
X_3853_ _0695_ VPWR _0700_ VGND _0696_ _0698_ sg13g2_o21ai_1
X_3784_ _0634_ _0622_ _0632_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_280 VPWR VGND sg13g2_fill_1
X_5523_ net454 mac2.sum_lvl3_ff\[24\] _2261_ VPWR VGND sg13g2_xor2_1
X_5454_ VGND VPWR _2204_ _2206_ _2207_ _2205_ sg13g2_a21oi_1
X_5385_ net317 mac1.sum_lvl3_ff\[25\] _2154_ VPWR VGND sg13g2_xor2_1
X_4405_ _1232_ _1204_ _1231_ VPWR VGND sg13g2_nand2_1
X_4336_ _1127_ VPWR _1164_ VGND _1085_ _1128_ sg13g2_o21ai_1
X_4267_ net817 net814 net858 net857 _1097_ VPWR VGND sg13g2_and4_1
X_3218_ _2809_ _2778_ _2807_ VPWR VGND sg13g2_xnor2_1
X_6006_ net1085 VGND VPWR _0111_ mac1.products_ff\[15\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_4198_ _1030_ net812 net866 VPWR VGND sg13g2_nand2_1
XFILLER_39_151 VPWR VGND sg13g2_fill_1
X_3149_ _2741_ _2733_ _2739_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_379 VPWR VGND sg13g2_decap_4
XFILLER_3_935 VPWR VGND sg13g2_decap_8
XFILLER_46_1001 VPWR VGND sg13g2_decap_8
Xhold280 mac2.sum_lvl2_ff\[2\] VPWR VGND net320 sg13g2_dlygate4sd3_1
XFILLER_49_64 VPWR VGND sg13g2_fill_1
Xhold291 DP_4.matrix\[38\] VPWR VGND net331 sg13g2_dlygate4sd3_1
XFILLER_49_97 VPWR VGND sg13g2_fill_2
Xfanout760 net762 net760 VPWR VGND sg13g2_buf_8
Xfanout782 net309 net782 VPWR VGND sg13g2_buf_8
Xfanout793 net795 net793 VPWR VGND sg13g2_buf_2
Xfanout771 net772 net771 VPWR VGND sg13g2_buf_8
XFILLER_10_780 VPWR VGND sg13g2_fill_2
XFILLER_46_4 VPWR VGND sg13g2_fill_1
X_5170_ _1964_ _1953_ _1965_ VPWR VGND sg13g2_xor2_1
X_4121_ _0960_ net907 net1009 VPWR VGND sg13g2_nand2_1
X_4052_ _0894_ _0874_ _0893_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_600 VPWR VGND sg13g2_decap_8
X_3003_ _2601_ _2594_ _2600_ VPWR VGND sg13g2_nand2_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_36_143 VPWR VGND sg13g2_fill_1
XFILLER_25_828 VPWR VGND sg13g2_fill_2
X_4954_ _1753_ _1752_ _1755_ VPWR VGND sg13g2_xor2_1
X_3905_ _0751_ _0749_ _0750_ VPWR VGND sg13g2_nand2_1
XFILLER_20_500 VPWR VGND sg13g2_fill_1
X_4885_ _1681_ _1683_ _1692_ VPWR VGND sg13g2_and2_1
X_3836_ _0660_ VPWR _0683_ VGND _0637_ _0658_ sg13g2_o21ai_1
X_3767_ _0618_ net973 net924 net918 net975 VPWR VGND sg13g2_a22oi_1
X_5506_ _0038_ _2247_ net532 VPWR VGND sg13g2_xnor2_1
X_6486_ net1018 VGND VPWR net349 mac2.total_sum\[14\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_3698_ _0554_ _0553_ _0555_ VPWR VGND sg13g2_nor2b_1
X_5437_ _2194_ net291 net267 VPWR VGND sg13g2_nand2_1
X_5368_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] _2141_ VPWR VGND sg13g2_nor2_1
XFILLER_0_927 VPWR VGND sg13g2_decap_8
X_5299_ _0007_ _2084_ net333 VPWR VGND sg13g2_xnor2_1
X_4319_ _1137_ _1145_ _1147_ _1148_ VPWR VGND sg13g2_or3_1
XFILLER_42_168 VPWR VGND sg13g2_fill_2
XFILLER_11_566 VPWR VGND sg13g2_fill_1
XFILLER_11_588 VPWR VGND sg13g2_fill_2
XFILLER_3_743 VPWR VGND sg13g2_fill_2
XFILLER_39_909 VPWR VGND sg13g2_decap_8
XFILLER_47_953 VPWR VGND sg13g2_decap_8
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_33_102 VPWR VGND sg13g2_fill_2
X_4670_ _1445_ VPWR _1484_ VGND _1446_ _1447_ sg13g2_o21ai_1
X_3621_ _0479_ _0475_ _0480_ VPWR VGND sg13g2_xor2_1
X_3552_ VGND VPWR _0409_ _0410_ _0413_ _0404_ sg13g2_a21oi_1
X_6340_ net1055 VGND VPWR _0085_ mac2.products_ff\[1\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3483_ _0345_ _0344_ _0112_ VPWR VGND sg13g2_xor2_1
X_6271_ net1033 VGND VPWR net97 mac2.sum_lvl1_ff\[84\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_5222_ _2015_ net841 net783 VPWR VGND sg13g2_nand2_1
X_5153_ VGND VPWR _1948_ _1946_ _1906_ sg13g2_or2_1
X_4104_ _0903_ _0943_ _0944_ VPWR VGND sg13g2_nor2_1
XFILLER_38_942 VPWR VGND sg13g2_decap_8
X_5084_ _1881_ _1874_ _1879_ _1880_ VPWR VGND sg13g2_and3_1
X_4035_ _0877_ net915 net1008 VPWR VGND sg13g2_nand2_1
XFILLER_36_1011 VPWR VGND sg13g2_decap_8
X_5986_ net1033 VGND VPWR net9 DP_3.Q_range.out_data\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_4937_ _1738_ net787 net854 net789 net852 VPWR VGND sg13g2_a22oi_1
X_4868_ _1638_ _1675_ _1676_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_341 VPWR VGND sg13g2_fill_2
X_3819_ _0663_ _0664_ _0666_ _0667_ VPWR VGND sg13g2_or3_1
X_4799_ _1592_ _1585_ _1553_ _1609_ VPWR VGND sg13g2_a21o_2
X_6469_ net1028 VGND VPWR net513 mac2.sum_lvl3_ff\[13\] clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_43_1004 VPWR VGND sg13g2_decap_8
XFILLER_0_724 VPWR VGND sg13g2_fill_1
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_47_227 VPWR VGND sg13g2_fill_2
XFILLER_16_614 VPWR VGND sg13g2_fill_1
XFILLER_16_625 VPWR VGND sg13g2_fill_1
XFILLER_29_986 VPWR VGND sg13g2_decap_8
XFILLER_44_956 VPWR VGND sg13g2_decap_8
XFILLER_8_879 VPWR VGND sg13g2_fill_1
XFILLER_3_562 VPWR VGND sg13g2_fill_1
XFILLER_3_551 VPWR VGND sg13g2_fill_2
XFILLER_38_227 VPWR VGND sg13g2_fill_2
XFILLER_47_772 VPWR VGND sg13g2_decap_4
XFILLER_35_901 VPWR VGND sg13g2_decap_8
XFILLER_34_411 VPWR VGND sg13g2_fill_2
X_5840_ VGND VPWR net756 _2539_ _0177_ _2538_ sg13g2_a21oi_1
XFILLER_35_978 VPWR VGND sg13g2_decap_8
X_5771_ _2478_ _2458_ _2477_ VPWR VGND sg13g2_nand2b_1
X_2983_ VPWR _2587_ DP_3.I_range.out_data\[3\] VGND sg13g2_inv_1
X_4722_ VGND VPWR _1534_ _1502_ _1500_ sg13g2_or2_1
X_4653_ _1463_ _1464_ _1466_ _1467_ VPWR VGND sg13g2_or3_1
X_3604_ _0464_ _0430_ _0463_ VPWR VGND sg13g2_nand2b_1
X_4584_ _1400_ net876 net835 net879 net832 VPWR VGND sg13g2_a22oi_1
X_6323_ net1012 VGND VPWR net284 mac1.total_sum\[0\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3535_ _0369_ VPWR _0396_ VGND _0360_ _0370_ sg13g2_o21ai_1
X_3466_ net933 net983 net938 _0329_ VPWR VGND net981 sg13g2_nand4_1
X_6254_ net1019 VGND VPWR net176 mac1.sum_lvl1_ff\[83\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5205_ _1999_ _1977_ _1998_ VPWR VGND sg13g2_xnor2_1
X_6185_ net1069 VGND VPWR net162 mac1.sum_lvl2_ff\[6\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3397_ _2978_ _2977_ _2970_ VPWR VGND sg13g2_nand2b_1
X_5136_ _1932_ _1901_ _1931_ VPWR VGND sg13g2_nand2_1
X_5067_ _1864_ _1856_ _1862_ VPWR VGND sg13g2_xnor2_1
X_4018_ _0859_ _0850_ _0861_ VPWR VGND sg13g2_xor2_1
XFILLER_26_901 VPWR VGND sg13g2_decap_8
XFILLER_38_783 VPWR VGND sg13g2_fill_2
XFILLER_26_978 VPWR VGND sg13g2_decap_8
X_5969_ net840 _0243_ VPWR VGND sg13g2_buf_1
XFILLER_41_948 VPWR VGND sg13g2_decap_8
XFILLER_32_12 VPWR VGND sg13g2_fill_2
XFILLER_40_469 VPWR VGND sg13g2_decap_4
XFILLER_21_650 VPWR VGND sg13g2_decap_8
XFILLER_0_543 VPWR VGND sg13g2_fill_2
XFILLER_17_989 VPWR VGND sg13g2_decap_8
XFILLER_32_948 VPWR VGND sg13g2_decap_8
XFILLER_8_676 VPWR VGND sg13g2_fill_2
Xhold109 mac1.products_ff\[77\] VPWR VGND net149 sg13g2_dlygate4sd3_1
X_3320_ _2851_ _2907_ _2908_ VPWR VGND sg13g2_nor2b_1
X_3251_ _2839_ _2830_ _2841_ VPWR VGND sg13g2_xor2_1
X_3182_ _2771_ _2770_ _2772_ _2774_ VPWR VGND sg13g2_a21o_1
XFILLER_14_2 VPWR VGND sg13g2_fill_1
X_5823_ VGND VPWR _2526_ _2527_ _0169_ _2528_ sg13g2_a21oi_1
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
X_5754_ net871 net886 net780 _2461_ VPWR VGND sg13g2_mux2_1
X_5685_ _2393_ _2390_ _2389_ _2394_ VPWR VGND sg13g2_a21o_1
X_4705_ _1515_ _1516_ _1497_ _1518_ VPWR VGND sg13g2_nand3_1
X_4636_ _1450_ net820 DP_3.matrix\[0\] net821 net885 VPWR VGND sg13g2_a22oi_1
XFILLER_2_808 VPWR VGND sg13g2_fill_1
X_6306_ net1082 VGND VPWR net287 mac1.sum_lvl3_ff\[15\] clknet_leaf_46_clk sg13g2_dfrbpq_2
X_4567_ _1383_ _1373_ _1384_ VPWR VGND sg13g2_xor2_1
X_3518_ _0377_ _0376_ _0346_ _0380_ VPWR VGND sg13g2_a21o_1
X_4498_ _1293_ _1319_ _1321_ VPWR VGND sg13g2_and2_1
X_3449_ _0313_ _0312_ _0311_ VPWR VGND sg13g2_nand2b_1
X_6237_ net1030 VGND VPWR net52 mac2.sum_lvl2_ff\[48\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6168_ net1068 VGND VPWR net177 mac1.sum_lvl1_ff\[41\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5119_ _1915_ net787 net841 VPWR VGND sg13g2_nand2_1
XFILLER_40_1018 VPWR VGND sg13g2_decap_8
X_6099_ net1047 VGND VPWR _0219_ DP_2.matrix\[79\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_49_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_27 VPWR VGND sg13g2_fill_2
XFILLER_1_885 VPWR VGND sg13g2_decap_8
XFILLER_36_517 VPWR VGND sg13g2_fill_2
XFILLER_9_952 VPWR VGND sg13g2_decap_8
X_5470_ VGND VPWR _2219_ _2220_ _2217_ net507 sg13g2_a21oi_2
X_4421_ _1246_ _1243_ _1247_ VPWR VGND sg13g2_xor2_1
X_4352_ VGND VPWR _1180_ _1179_ _1132_ sg13g2_or2_1
X_3303_ _2891_ net945 net889 VPWR VGND sg13g2_nand2_1
X_4283_ VGND VPWR _1110_ _1111_ _1113_ _1081_ sg13g2_a21oi_1
X_3234_ VGND VPWR _2824_ _2822_ _2783_ sg13g2_or2_1
X_6022_ net1085 VGND VPWR _0122_ mac1.products_ff\[83\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_39_333 VPWR VGND sg13g2_fill_2
X_3165_ _2752_ VPWR _2757_ VGND _2753_ _2755_ sg13g2_o21ai_1
X_3096_ _2690_ _2666_ _2689_ VPWR VGND sg13g2_xnor2_1
X_5806_ net808 net779 _2512_ VPWR VGND sg13g2_nor2_1
X_3998_ _0841_ net974 net1004 VPWR VGND sg13g2_nand2_1
X_5737_ VGND VPWR _2442_ _2443_ _0163_ _2444_ sg13g2_a21oi_1
X_5668_ net983 DP_1.matrix\[41\] net775 _2377_ VPWR VGND sg13g2_mux2_1
X_5599_ net30 _2317_ _2319_ VPWR VGND sg13g2_xnor2_1
X_4619_ _1429_ VPWR _1434_ VGND _1430_ _1432_ sg13g2_o21ai_1
Xhold451 DP_1.matrix\[39\] VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold462 DP_1.matrix\[6\] VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold440 _2131_ VPWR VGND net480 sg13g2_dlygate4sd3_1
Xhold495 mac1.sum_lvl2_ff\[12\] VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold484 mac2.sum_lvl2_ff\[6\] VPWR VGND net524 sg13g2_dlygate4sd3_1
Xhold473 _0036_ VPWR VGND net513 sg13g2_dlygate4sd3_1
Xfanout931 DP_2.matrix\[2\] net931 VPWR VGND sg13g2_buf_1
Xfanout920 net921 net920 VPWR VGND sg13g2_buf_1
Xfanout942 net943 net942 VPWR VGND sg13g2_buf_1
Xfanout986 net510 net986 VPWR VGND sg13g2_buf_8
Xfanout953 net326 net953 VPWR VGND sg13g2_buf_8
Xfanout975 net412 net975 VPWR VGND sg13g2_buf_8
Xfanout964 net965 net964 VPWR VGND sg13g2_buf_1
Xfanout997 net316 net997 VPWR VGND sg13g2_buf_8
XFILLER_13_200 VPWR VGND sg13g2_fill_1
XFILLER_41_542 VPWR VGND sg13g2_fill_1
XFILLER_41_575 VPWR VGND sg13g2_decap_4
XFILLER_9_237 VPWR VGND sg13g2_fill_2
XFILLER_13_299 VPWR VGND sg13g2_fill_1
XFILLER_6_933 VPWR VGND sg13g2_decap_8
XFILLER_5_410 VPWR VGND sg13g2_fill_1
Xclkload18 clknet_leaf_57_clk clkload18/Y VPWR VGND sg13g2_inv_4
XFILLER_5_465 VPWR VGND sg13g2_fill_1
XFILLER_49_642 VPWR VGND sg13g2_decap_8
XFILLER_0_170 VPWR VGND sg13g2_fill_2
XFILLER_45_881 VPWR VGND sg13g2_decap_8
X_4970_ _1765_ VPWR _1770_ VGND _1766_ _1768_ sg13g2_o21ai_1
XFILLER_44_391 VPWR VGND sg13g2_fill_2
X_3921_ net914 net968 net912 net966 _0766_ VPWR VGND sg13g2_and4_1
X_3852_ _0695_ _0696_ _0698_ _0699_ VPWR VGND sg13g2_or3_1
XFILLER_32_586 VPWR VGND sg13g2_fill_1
X_3783_ _0633_ _0632_ _0622_ VPWR VGND sg13g2_nand2b_1
X_5522_ mac2.sum_lvl3_ff\[24\] mac2.sum_lvl3_ff\[4\] _2260_ VPWR VGND sg13g2_and2_1
X_5453_ net462 _2204_ _0042_ VPWR VGND sg13g2_xor2_1
X_5384_ mac1.sum_lvl3_ff\[25\] net317 _2153_ VPWR VGND sg13g2_nor2_1
X_4404_ _1229_ _1205_ _1231_ VPWR VGND sg13g2_xor2_1
X_4335_ _0136_ _1118_ _1162_ VPWR VGND sg13g2_xnor2_1
X_4266_ _1096_ net812 net861 VPWR VGND sg13g2_nand2_1
X_3217_ _2808_ _2778_ _2807_ VPWR VGND sg13g2_nand2_1
X_6005_ net1085 VGND VPWR _0110_ mac1.products_ff\[14\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_4197_ _1010_ VPWR _1029_ VGND _1008_ _1011_ sg13g2_o21ai_1
X_3148_ _2740_ _2733_ _2739_ VPWR VGND sg13g2_nand2_1
X_3079_ _2673_ _2668_ _2671_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_892 VPWR VGND sg13g2_decap_8
XFILLER_40_45 VPWR VGND sg13g2_decap_8
XFILLER_3_914 VPWR VGND sg13g2_decap_8
Xhold270 DP_2.matrix\[74\] VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold292 mac1.sum_lvl2_ff\[1\] VPWR VGND net332 sg13g2_dlygate4sd3_1
Xhold281 _2200_ VPWR VGND net321 sg13g2_dlygate4sd3_1
XFILLER_49_76 VPWR VGND sg13g2_decap_8
XFILLER_46_601 VPWR VGND sg13g2_fill_2
Xfanout761 net762 net761 VPWR VGND sg13g2_buf_8
Xfanout794 net796 net794 VPWR VGND sg13g2_buf_1
Xfanout783 net784 net783 VPWR VGND sg13g2_buf_8
Xfanout772 _2372_ net772 VPWR VGND sg13g2_buf_8
XFILLER_46_634 VPWR VGND sg13g2_fill_1
XFILLER_18_347 VPWR VGND sg13g2_fill_1
XFILLER_45_199 VPWR VGND sg13g2_fill_2
XFILLER_14_597 VPWR VGND sg13g2_fill_1
XFILLER_6_741 VPWR VGND sg13g2_fill_2
X_4120_ _0959_ net964 DP_2.matrix\[44\] VPWR VGND sg13g2_nand2_1
X_4051_ _0891_ _0881_ _0893_ VPWR VGND sg13g2_xor2_1
X_3002_ _2599_ _2596_ _2600_ VPWR VGND sg13g2_xor2_1
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_37_667 VPWR VGND sg13g2_fill_2
X_4953_ _1754_ _1752_ _1753_ VPWR VGND sg13g2_nand2_1
XFILLER_36_199 VPWR VGND sg13g2_fill_2
X_3904_ _0711_ VPWR _0750_ VGND _0712_ _0713_ sg13g2_o21ai_1
X_4884_ _1689_ _1665_ _1690_ _1691_ VPWR VGND sg13g2_a21o_1
XFILLER_32_383 VPWR VGND sg13g2_fill_1
XFILLER_33_895 VPWR VGND sg13g2_decap_8
X_3835_ _0682_ _0674_ _0678_ VPWR VGND sg13g2_nand2_1
X_3766_ net924 net975 net918 net973 _0617_ VPWR VGND sg13g2_and4_1
X_5505_ _2248_ mac2.sum_lvl2_ff\[34\] net531 VPWR VGND sg13g2_xnor2_1
X_6485_ net1018 VGND VPWR net401 mac2.total_sum\[13\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5436_ net283 mac1.sum_lvl3_ff\[20\] _0016_ VPWR VGND sg13g2_xor2_1
X_3697_ VGND VPWR _0508_ _0513_ _0554_ _0527_ sg13g2_a21oi_1
X_5367_ _2140_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_0_906 VPWR VGND sg13g2_decap_8
X_5298_ net332 mac1.sum_lvl2_ff\[20\] _2087_ VPWR VGND sg13g2_xor2_1
X_4318_ VGND VPWR _1143_ _1144_ _1147_ _1138_ sg13g2_a21oi_1
XFILLER_47_409 VPWR VGND sg13g2_fill_1
X_4249_ VGND VPWR _1021_ _1047_ _1080_ _1046_ sg13g2_a21oi_1
XFILLER_3_777 VPWR VGND sg13g2_fill_1
XFILLER_2_254 VPWR VGND sg13g2_fill_2
XFILLER_47_932 VPWR VGND sg13g2_decap_8
XFILLER_20_1005 VPWR VGND sg13g2_decap_8
XFILLER_15_895 VPWR VGND sg13g2_fill_2
X_3620_ _0479_ _0435_ _0477_ VPWR VGND sg13g2_xnor2_1
X_3551_ _0409_ _0410_ _0404_ _0412_ VPWR VGND sg13g2_nand3_1
X_3482_ VGND VPWR _0286_ _0312_ _0345_ _0311_ sg13g2_a21oi_1
X_6270_ net1026 VGND VPWR net209 mac2.sum_lvl1_ff\[83\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5221_ _2014_ net841 net781 VPWR VGND sg13g2_nand2_1
X_5152_ _1947_ net846 net783 VPWR VGND sg13g2_nand2_1
X_4103_ _0943_ _0934_ _0942_ VPWR VGND sg13g2_xnor2_1
X_5083_ _1875_ VPWR _1880_ VGND _1876_ _1878_ sg13g2_o21ai_1
XFILLER_38_921 VPWR VGND sg13g2_decap_8
X_4034_ _0876_ net910 net964 VPWR VGND sg13g2_nand2_1
XFILLER_38_998 VPWR VGND sg13g2_decap_8
X_5985_ net782 _0267_ VPWR VGND sg13g2_buf_1
XFILLER_21_821 VPWR VGND sg13g2_fill_2
X_4936_ _0092_ _1723_ _1736_ VPWR VGND sg13g2_xnor2_1
X_4867_ _1675_ _1670_ _1673_ VPWR VGND sg13g2_xnor2_1
X_3818_ _0666_ net967 net923 net969 net921 VPWR VGND sg13g2_a22oi_1
X_4798_ _1594_ VPWR _1608_ VGND _1583_ _1595_ sg13g2_o21ai_1
X_3749_ _0602_ _0589_ _0604_ VPWR VGND sg13g2_xor2_1
X_6468_ net1029 VGND VPWR _0035_ mac2.sum_lvl3_ff\[12\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6399_ net1093 VGND VPWR net263 mac2.sum_lvl1_ff\[12\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_5419_ _2181_ mac1.sum_lvl3_ff\[32\] net323 VPWR VGND sg13g2_nand2_1
XFILLER_29_965 VPWR VGND sg13g2_decap_8
XFILLER_44_935 VPWR VGND sg13g2_decap_8
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_1010 VPWR VGND sg13g2_decap_8
XFILLER_35_957 VPWR VGND sg13g2_decap_8
XFILLER_43_990 VPWR VGND sg13g2_decap_8
X_5770_ _2477_ _2476_ _2472_ VPWR VGND sg13g2_nand2b_1
XFILLER_34_478 VPWR VGND sg13g2_fill_2
X_4721_ _1492_ VPWR _1533_ VGND _1451_ _1490_ sg13g2_o21ai_1
X_4652_ _1466_ net873 net836 net874 net831 VPWR VGND sg13g2_a22oi_1
X_3603_ _0463_ _0431_ _0461_ VPWR VGND sg13g2_xnor2_1
X_4583_ net832 net878 net835 _1399_ VPWR VGND net876 sg13g2_nand4_1
X_6322_ net1034 VGND VPWR net174 mac2.sum_lvl3_ff\[35\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3534_ _0395_ _0350_ _0394_ VPWR VGND sg13g2_xnor2_1
X_3465_ net938 net935 net983 net981 _0328_ VPWR VGND sg13g2_and4_1
X_6253_ net1019 VGND VPWR net225 mac1.sum_lvl1_ff\[82\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5204_ _1996_ _1984_ _1998_ VPWR VGND sg13g2_xor2_1
X_3396_ _2975_ _2976_ _2977_ VPWR VGND sg13g2_nor2b_1
X_6184_ net1068 VGND VPWR net157 mac1.sum_lvl2_ff\[5\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5135_ _1930_ _1912_ _1931_ VPWR VGND sg13g2_xor2_1
X_5066_ _1863_ _1856_ _1862_ VPWR VGND sg13g2_nand2_1
X_4017_ _0860_ _0850_ _0859_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_957 VPWR VGND sg13g2_decap_8
XFILLER_25_445 VPWR VGND sg13g2_fill_1
X_5968_ net843 _0242_ VPWR VGND sg13g2_buf_1
XFILLER_41_927 VPWR VGND sg13g2_decap_8
X_4919_ _1721_ _1718_ _1722_ VPWR VGND sg13g2_xor2_1
X_5899_ _2509_ _2499_ _2577_ VPWR VGND sg13g2_xor2_1
XFILLER_4_338 VPWR VGND sg13g2_fill_1
XFILLER_29_740 VPWR VGND sg13g2_fill_1
XFILLER_17_913 VPWR VGND sg13g2_decap_8
XFILLER_16_412 VPWR VGND sg13g2_fill_1
XFILLER_17_968 VPWR VGND sg13g2_decap_8
XFILLER_44_787 VPWR VGND sg13g2_fill_2
XFILLER_32_927 VPWR VGND sg13g2_decap_8
XFILLER_4_883 VPWR VGND sg13g2_fill_2
X_3250_ _2840_ _2830_ _2839_ VPWR VGND sg13g2_nand2b_1
X_3181_ _2771_ _2772_ _2770_ _2773_ VPWR VGND sg13g2_nand3_1
XFILLER_39_504 VPWR VGND sg13g2_fill_2
XFILLER_35_732 VPWR VGND sg13g2_decap_4
X_5822_ _2493_ _2527_ _2528_ VPWR VGND sg13g2_nor2_1
XFILLER_35_798 VPWR VGND sg13g2_decap_4
X_5753_ _2460_ _2459_ net769 net765 net421 VPWR VGND sg13g2_a22oi_1
X_4704_ _1517_ _1497_ _1515_ _1516_ VPWR VGND sg13g2_and3_1
X_5684_ _2392_ VPWR _2393_ VGND net989 net776 sg13g2_o21ai_1
X_4635_ _1426_ VPWR _1449_ VGND _1391_ _1424_ sg13g2_o21ai_1
X_4566_ _1383_ _1381_ _1382_ VPWR VGND sg13g2_nand2_1
X_3517_ VGND VPWR _0376_ _0377_ _0379_ _0346_ sg13g2_a21oi_1
X_6305_ net1047 VGND VPWR net470 mac1.sum_lvl3_ff\[14\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_4497_ _1320_ _1319_ _0131_ VPWR VGND sg13g2_xor2_1
X_3448_ _0284_ VPWR _0312_ VGND _0308_ _0309_ sg13g2_o21ai_1
X_6236_ net1028 VGND VPWR net42 mac2.sum_lvl2_ff\[47\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3379_ _2962_ net932 net993 net991 net937 VPWR VGND sg13g2_a22oi_1
X_6167_ net1068 VGND VPWR net86 mac1.sum_lvl1_ff\[40\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5118_ _1914_ net846 net785 VPWR VGND sg13g2_nand2_1
X_6098_ net1048 VGND VPWR _0218_ DP_2.matrix\[78\] clknet_leaf_60_clk sg13g2_dfrbpq_2
XFILLER_26_710 VPWR VGND sg13g2_decap_4
X_5049_ _1823_ VPWR _1847_ VGND _1843_ _1845_ sg13g2_o21ai_1
XFILLER_43_67 VPWR VGND sg13g2_fill_1
XFILLER_41_779 VPWR VGND sg13g2_fill_2
XFILLER_5_614 VPWR VGND sg13g2_decap_4
XFILLER_44_540 VPWR VGND sg13g2_decap_4
XFILLER_16_242 VPWR VGND sg13g2_fill_2
XFILLER_44_584 VPWR VGND sg13g2_decap_8
XFILLER_44_595 VPWR VGND sg13g2_fill_2
XFILLER_9_931 VPWR VGND sg13g2_decap_8
XFILLER_13_982 VPWR VGND sg13g2_decap_8
X_4420_ _1246_ _1220_ _1244_ VPWR VGND sg13g2_xnor2_1
X_4351_ _1179_ net809 net858 VPWR VGND sg13g2_nand2_1
X_3302_ _2890_ net945 net887 VPWR VGND sg13g2_nand2_1
X_4282_ _1110_ _1111_ _1081_ _1112_ VPWR VGND sg13g2_nand3_1
X_3233_ _2823_ net950 net889 VPWR VGND sg13g2_nand2_1
X_6021_ net1083 VGND VPWR _0121_ mac1.products_ff\[82\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_3164_ _2752_ _2753_ _2755_ _2756_ VPWR VGND sg13g2_or3_1
XFILLER_12_0 VPWR VGND sg13g2_fill_2
X_3095_ _2689_ _2686_ _2688_ VPWR VGND sg13g2_nand2_1
XFILLER_35_540 VPWR VGND sg13g2_decap_4
XFILLER_23_713 VPWR VGND sg13g2_decap_4
X_5805_ _2511_ net788 net766 VPWR VGND sg13g2_nand2_1
X_3997_ _0813_ VPWR _0840_ VGND _0811_ _0814_ sg13g2_o21ai_1
XFILLER_11_908 VPWR VGND sg13g2_decap_4
X_5736_ _2411_ _2443_ _2444_ VPWR VGND sg13g2_nor2_1
X_5667_ _2590_ _2375_ net756 _2376_ VPWR VGND sg13g2_mux2_1
X_4618_ _1429_ _1430_ _1432_ _1433_ VPWR VGND sg13g2_or3_1
X_5598_ mac2.total_sum\[5\] mac1.total_sum\[5\] _2319_ VPWR VGND sg13g2_xor2_1
Xhold452 DP_3.matrix\[40\] VPWR VGND net492 sg13g2_dlygate4sd3_1
Xhold463 DP_1.matrix\[5\] VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold441 _0004_ VPWR VGND net481 sg13g2_dlygate4sd3_1
Xhold430 _0005_ VPWR VGND net470 sg13g2_dlygate4sd3_1
X_4549_ _1367_ _1366_ _1356_ VPWR VGND sg13g2_nand2b_1
Xhold474 mac1.sum_lvl2_ff\[6\] VPWR VGND net514 sg13g2_dlygate4sd3_1
Xhold496 _2128_ VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold485 _2211_ VPWR VGND net525 sg13g2_dlygate4sd3_1
Xfanout932 net936 net932 VPWR VGND sg13g2_buf_8
Xfanout921 DP_2.matrix\[37\] net921 VPWR VGND sg13g2_buf_1
Xfanout943 DP_1.matrix\[79\] net943 VPWR VGND sg13g2_buf_1
X_6219_ net1014 VGND VPWR net216 mac1.sum_lvl2_ff\[46\] clknet_leaf_2_clk sg13g2_dfrbpq_1
Xfanout910 net911 net910 VPWR VGND sg13g2_buf_8
Xfanout976 net412 net976 VPWR VGND sg13g2_buf_1
Xfanout954 net955 net954 VPWR VGND sg13g2_buf_8
Xfanout965 net528 net965 VPWR VGND sg13g2_buf_2
Xfanout998 DP_3.matrix\[80\] net998 VPWR VGND sg13g2_buf_1
Xfanout987 net988 net987 VPWR VGND sg13g2_buf_8
XFILLER_13_245 VPWR VGND sg13g2_fill_1
XFILLER_10_985 VPWR VGND sg13g2_decap_8
Xclkload19 clkload19/Y clknet_leaf_59_clk VPWR VGND sg13g2_inv_2
XFILLER_6_989 VPWR VGND sg13g2_decap_8
XFILLER_49_621 VPWR VGND sg13g2_decap_8
XFILLER_0_193 VPWR VGND sg13g2_decap_4
XFILLER_0_182 VPWR VGND sg13g2_fill_1
XFILLER_48_186 VPWR VGND sg13g2_fill_2
X_3920_ _0765_ net912 net967 VPWR VGND sg13g2_nand2_1
X_3851_ _0698_ net965 net922 net967 net920 VPWR VGND sg13g2_a22oi_1
X_3782_ _0632_ _0623_ _0630_ VPWR VGND sg13g2_xnor2_1
X_5521_ _2257_ VPWR _2259_ VGND _2256_ _2258_ sg13g2_o21ai_1
XFILLER_30_1018 VPWR VGND sg13g2_decap_8
X_5452_ net461 mac2.sum_lvl2_ff\[23\] _2206_ VPWR VGND sg13g2_xor2_1
X_5383_ VGND VPWR _2149_ _2151_ _2152_ _2150_ sg13g2_a21oi_1
X_4403_ _1230_ _1205_ _1229_ VPWR VGND sg13g2_nand2_1
X_4334_ _1117_ _1162_ _1116_ _1163_ VPWR VGND sg13g2_nand3_1
XFILLER_8_1008 VPWR VGND sg13g2_decap_8
X_6004_ net1082 VGND VPWR _0109_ mac1.products_ff\[13\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_4265_ _1064_ VPWR _1095_ VGND _1062_ _1065_ sg13g2_o21ai_1
X_3216_ _2806_ _2789_ _2807_ VPWR VGND sg13g2_xor2_1
X_4196_ _1026_ _1023_ _1028_ VPWR VGND sg13g2_xor2_1
XFILLER_39_120 VPWR VGND sg13g2_fill_1
X_3147_ _2739_ _2734_ _2737_ VPWR VGND sg13g2_xnor2_1
X_3078_ _2672_ _2671_ _2668_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_871 VPWR VGND sg13g2_decap_8
XFILLER_39_1021 VPWR VGND sg13g2_decap_8
XFILLER_24_36 VPWR VGND sg13g2_fill_1
X_5719_ VPWR _2427_ _2426_ VGND sg13g2_inv_1
XFILLER_40_57 VPWR VGND sg13g2_fill_2
Xhold260 DP_4.matrix\[75\] VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold271 mac2.sum_lvl3_ff\[12\] VPWR VGND net311 sg13g2_dlygate4sd3_1
Xhold293 _2087_ VPWR VGND net333 sg13g2_dlygate4sd3_1
Xhold282 _0040_ VPWR VGND net322 sg13g2_dlygate4sd3_1
XFILLER_49_99 VPWR VGND sg13g2_fill_1
Xfanout784 net315 net784 VPWR VGND sg13g2_buf_2
Xfanout773 net774 net773 VPWR VGND sg13g2_buf_8
Xfanout762 _2487_ net762 VPWR VGND sg13g2_buf_8
XFILLER_45_101 VPWR VGND sg13g2_fill_1
Xfanout795 net796 net795 VPWR VGND sg13g2_buf_2
XFILLER_45_145 VPWR VGND sg13g2_fill_2
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_42_841 VPWR VGND sg13g2_fill_2
XFILLER_41_351 VPWR VGND sg13g2_fill_1
XFILLER_42_896 VPWR VGND sg13g2_decap_8
XFILLER_5_241 VPWR VGND sg13g2_fill_1
XFILLER_2_992 VPWR VGND sg13g2_decap_8
X_4050_ _0881_ _0891_ _0892_ VPWR VGND sg13g2_nor2_1
X_3001_ _2597_ _2598_ _2599_ VPWR VGND sg13g2_nor2_1
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
XFILLER_24_318 VPWR VGND sg13g2_decap_4
XFILLER_45_690 VPWR VGND sg13g2_fill_1
X_4952_ _1753_ _1733_ _1735_ VPWR VGND sg13g2_nand2_1
X_4883_ VGND VPWR _1660_ _1686_ _1690_ _1685_ sg13g2_a21oi_1
X_3903_ _0748_ _0685_ _0749_ VPWR VGND sg13g2_xor2_1
XFILLER_33_874 VPWR VGND sg13g2_decap_8
X_3834_ _0116_ _0654_ _0681_ VPWR VGND sg13g2_xnor2_1
X_3765_ net977 net916 _0616_ VPWR VGND sg13g2_and2_1
X_5504_ _2244_ VPWR _2247_ VGND _2243_ _2245_ sg13g2_o21ai_1
XFILLER_9_591 VPWR VGND sg13g2_decap_8
X_3696_ _0551_ _0540_ _0553_ VPWR VGND sg13g2_xor2_1
X_6484_ net1018 VGND VPWR net313 mac2.total_sum\[12\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_10_27 VPWR VGND sg13g2_fill_2
X_5435_ _0022_ _2192_ net410 VPWR VGND sg13g2_xnor2_1
X_5366_ _2139_ net429 net283 VPWR VGND sg13g2_nand2_1
X_5297_ mac1.sum_lvl2_ff\[20\] net332 _2086_ VPWR VGND sg13g2_nor2_1
X_4317_ _1143_ _1144_ _1138_ _1146_ VPWR VGND sg13g2_nand3_1
X_4248_ _1077_ _1049_ _1079_ VPWR VGND sg13g2_xor2_1
XFILLER_19_58 VPWR VGND sg13g2_fill_2
XFILLER_28_602 VPWR VGND sg13g2_fill_2
X_4179_ _1008_ _1009_ _1011_ _1012_ VPWR VGND sg13g2_or3_1
XFILLER_16_819 VPWR VGND sg13g2_fill_1
XFILLER_11_557 VPWR VGND sg13g2_decap_8
XFILLER_13_1024 VPWR VGND sg13g2_decap_4
XFILLER_2_211 VPWR VGND sg13g2_fill_1
XFILLER_47_911 VPWR VGND sg13g2_decap_8
XFILLER_46_421 VPWR VGND sg13g2_fill_2
XFILLER_19_646 VPWR VGND sg13g2_decap_4
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_988 VPWR VGND sg13g2_decap_8
XFILLER_14_340 VPWR VGND sg13g2_fill_1
XFILLER_25_90 VPWR VGND sg13g2_fill_1
XFILLER_41_181 VPWR VGND sg13g2_decap_8
XFILLER_30_899 VPWR VGND sg13g2_decap_8
X_3550_ _0411_ _0404_ _0409_ _0410_ VPWR VGND sg13g2_and3_1
X_5220_ _2013_ net846 net994 VPWR VGND sg13g2_nand2_1
X_3481_ _0342_ _0314_ _0344_ VPWR VGND sg13g2_xor2_1
X_5151_ _1946_ net846 net781 VPWR VGND sg13g2_nand2_1
X_5082_ _1875_ _1876_ _1878_ _1879_ VPWR VGND sg13g2_or3_1
X_4102_ _0942_ _0904_ _0940_ VPWR VGND sg13g2_xnor2_1
X_4033_ _0858_ _0851_ _0819_ _0875_ VPWR VGND sg13g2_a21o_1
XFILLER_38_900 VPWR VGND sg13g2_decap_8
XFILLER_38_977 VPWR VGND sg13g2_decap_8
XFILLER_24_104 VPWR VGND sg13g2_fill_2
X_5984_ net784 _0266_ VPWR VGND sg13g2_buf_1
X_4935_ _1723_ _1736_ _1737_ VPWR VGND sg13g2_nor2b_1
X_4866_ _1674_ _1673_ _1670_ VPWR VGND sg13g2_nand2b_1
X_4797_ _1580_ _1574_ _1582_ _1607_ VPWR VGND sg13g2_a21o_1
X_3817_ net921 net969 net923 _0665_ VPWR VGND net967 sg13g2_nand4_1
XFILLER_20_343 VPWR VGND sg13g2_fill_1
X_3748_ VGND VPWR _0603_ _0602_ _0589_ sg13g2_or2_1
XFILLER_4_509 VPWR VGND sg13g2_fill_2
X_3679_ _0524_ VPWR _0536_ VGND _0516_ _0525_ sg13g2_o21ai_1
X_6467_ net1028 VGND VPWR _0034_ mac2.sum_lvl3_ff\[11\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5418_ VPWR VGND _2178_ _2179_ _2171_ mac1.sum_lvl3_ff\[31\] _2180_ mac1.sum_lvl3_ff\[11\]
+ sg13g2_a221oi_1
X_6398_ net1090 VGND VPWR net93 mac2.sum_lvl1_ff\[11\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_5349_ _2127_ mac1.sum_lvl2_ff\[31\] mac1.sum_lvl2_ff\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_47_229 VPWR VGND sg13g2_fill_1
XFILLER_29_944 VPWR VGND sg13g2_decap_8
XFILLER_46_67 VPWR VGND sg13g2_fill_2
XFILLER_44_914 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_50_clk clknet_4_10_0_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
XFILLER_38_229 VPWR VGND sg13g2_fill_1
XFILLER_34_413 VPWR VGND sg13g2_fill_1
XFILLER_34_424 VPWR VGND sg13g2_fill_1
XFILLER_35_936 VPWR VGND sg13g2_decap_8
XFILLER_15_671 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_41_clk clknet_4_13_0_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4720_ _1518_ VPWR _1532_ VGND _1496_ _1519_ sg13g2_o21ai_1
X_4651_ net831 net874 net835 _1465_ VPWR VGND net873 sg13g2_nand4_1
X_3602_ _0462_ _0431_ _0461_ VPWR VGND sg13g2_nand2_1
X_4582_ net835 net832 net878 net876 _1398_ VPWR VGND sg13g2_and4_1
X_3533_ _0394_ _0386_ _0392_ VPWR VGND sg13g2_xnor2_1
X_6321_ net1034 VGND VPWR net241 mac2.sum_lvl3_ff\[34\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3464_ _0327_ net931 net986 VPWR VGND sg13g2_nand2_1
X_6252_ net1019 VGND VPWR net259 mac1.sum_lvl1_ff\[81\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5203_ _1984_ _1996_ _1997_ VPWR VGND sg13g2_nor2_1
X_6183_ net1068 VGND VPWR net101 mac1.sum_lvl2_ff\[4\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3395_ _2971_ VPWR _2976_ VGND _2972_ _2974_ sg13g2_o21ai_1
X_5134_ _1930_ _1913_ _1928_ VPWR VGND sg13g2_xnor2_1
X_5065_ _1862_ _1857_ _1860_ VPWR VGND sg13g2_xnor2_1
X_4016_ _0859_ _0851_ _0858_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_936 VPWR VGND sg13g2_decap_8
XFILLER_38_785 VPWR VGND sg13g2_fill_1
XFILLER_41_906 VPWR VGND sg13g2_decap_8
X_5967_ net274 _0241_ VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_32_clk clknet_4_13_0_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
X_4918_ _1719_ _1720_ _1721_ VPWR VGND sg13g2_nor2_1
XFILLER_32_14 VPWR VGND sg13g2_fill_1
X_5898_ _2576_ VPWR _0246_ VGND net759 _2575_ sg13g2_o21ai_1
X_4849_ _1658_ _1635_ _1657_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_947 VPWR VGND sg13g2_decap_8
XFILLER_44_766 VPWR VGND sg13g2_fill_1
XFILLER_32_906 VPWR VGND sg13g2_decap_8
XFILLER_25_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_4_5_0_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_31_427 VPWR VGND sg13g2_fill_2
XFILLER_31_449 VPWR VGND sg13g2_fill_1
XFILLER_12_652 VPWR VGND sg13g2_decap_8
XFILLER_11_162 VPWR VGND sg13g2_fill_1
XFILLER_40_983 VPWR VGND sg13g2_decap_8
XFILLER_22_80 VPWR VGND sg13g2_fill_2
XFILLER_22_91 VPWR VGND sg13g2_fill_2
X_3180_ _2725_ VPWR _2772_ VGND _2665_ _2726_ sg13g2_o21ai_1
X_5821_ _2527_ _2524_ net762 VPWR VGND sg13g2_nand2b_1
XFILLER_16_991 VPWR VGND sg13g2_decap_8
X_5752_ net865 net880 net780 _2459_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_14_clk clknet_4_6_0_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_4703_ _1504_ VPWR _1516_ VGND _1512_ _1514_ sg13g2_o21ai_1
X_5683_ VPWR _2392_ _2391_ VGND sg13g2_inv_1
XFILLER_31_983 VPWR VGND sg13g2_decap_8
X_4634_ _1440_ VPWR _1448_ VGND _1420_ _1441_ sg13g2_o21ai_1
X_4565_ _1380_ _1379_ _1374_ _1382_ VPWR VGND sg13g2_a21o_1
X_3516_ _0376_ _0377_ _0346_ _0378_ VPWR VGND sg13g2_nand3_1
X_6304_ net1042 VGND VPWR net481 mac1.sum_lvl3_ff\[13\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4496_ _1320_ _1292_ _1298_ VPWR VGND sg13g2_nand2_1
X_3447_ _0284_ _0308_ _0309_ _0311_ VPWR VGND sg13g2_nor3_1
X_6235_ net1028 VGND VPWR net104 mac2.sum_lvl2_ff\[46\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6166_ net1067 VGND VPWR net134 mac1.sum_lvl1_ff\[39\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3378_ _2961_ net991 net932 _0069_ VPWR VGND sg13g2_and3_2
X_6097_ net1043 VGND VPWR net89 mac1.sum_lvl1_ff\[0\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_5117_ _1882_ VPWR _1913_ VGND _1873_ _1883_ sg13g2_o21ai_1
X_5048_ _1823_ _1843_ _1845_ _1846_ VPWR VGND sg13g2_or3_1
XFILLER_14_906 VPWR VGND sg13g2_fill_1
XFILLER_26_744 VPWR VGND sg13g2_fill_2
XFILLER_41_725 VPWR VGND sg13g2_fill_2
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_41_769 VPWR VGND sg13g2_fill_2
XFILLER_22_983 VPWR VGND sg13g2_decap_8
XFILLER_49_825 VPWR VGND sg13g2_fill_2
XFILLER_48_335 VPWR VGND sg13g2_fill_2
XFILLER_36_508 VPWR VGND sg13g2_decap_4
XFILLER_1_1025 VPWR VGND sg13g2_decap_4
XFILLER_13_961 VPWR VGND sg13g2_decap_8
XFILLER_20_909 VPWR VGND sg13g2_decap_8
XFILLER_12_482 VPWR VGND sg13g2_decap_4
XFILLER_9_987 VPWR VGND sg13g2_decap_8
X_4350_ _1178_ net864 net806 VPWR VGND sg13g2_nand2_1
X_3301_ _2889_ net951 net1003 VPWR VGND sg13g2_nand2_1
X_4281_ _1088_ VPWR _1111_ VGND _1107_ _1109_ sg13g2_o21ai_1
X_3232_ _2822_ net949 net887 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_3_clk clknet_4_3_0_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_6020_ net1083 VGND VPWR _0120_ mac1.products_ff\[81\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_3163_ _2755_ net1006 net905 net941 net900 VPWR VGND sg13g2_a22oi_1
XFILLER_39_335 VPWR VGND sg13g2_fill_1
XFILLER_48_891 VPWR VGND sg13g2_decap_8
X_3094_ _2685_ _2684_ _2667_ _2688_ VPWR VGND sg13g2_a21o_1
X_5804_ _2510_ _2509_ _2499_ VPWR VGND sg13g2_nand2b_1
X_3996_ _0804_ VPWR _0839_ VGND _0801_ _0805_ sg13g2_o21ai_1
X_5735_ net756 VPWR _2443_ VGND _2439_ _2441_ sg13g2_o21ai_1
X_5666_ net764 net269 _2374_ _2375_ VPWR VGND sg13g2_a21o_1
X_4617_ _1432_ net874 net836 net876 net832 VPWR VGND sg13g2_a22oi_1
X_5597_ mac1.total_sum\[5\] mac2.total_sum\[5\] _2318_ VPWR VGND sg13g2_nor2_1
Xhold420 _0060_ VPWR VGND net460 sg13g2_dlygate4sd3_1
Xhold442 DP_4.matrix\[41\] VPWR VGND net482 sg13g2_dlygate4sd3_1
Xhold431 DP_2.matrix\[41\] VPWR VGND net471 sg13g2_dlygate4sd3_1
X_4548_ _1366_ _1357_ _1364_ VPWR VGND sg13g2_xnor2_1
Xhold453 DP_3.matrix\[3\] VPWR VGND net493 sg13g2_dlygate4sd3_1
X_4479_ _1303_ net856 net801 VPWR VGND sg13g2_nand2_1
Xhold464 DP_2.matrix\[39\] VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold475 _2101_ VPWR VGND net515 sg13g2_dlygate4sd3_1
Xfanout900 net901 net900 VPWR VGND sg13g2_buf_2
Xhold486 _2214_ VPWR VGND net526 sg13g2_dlygate4sd3_1
X_6218_ net1014 VGND VPWR net193 mac1.sum_lvl2_ff\[45\] clknet_leaf_1_clk sg13g2_dfrbpq_1
Xfanout922 net923 net922 VPWR VGND sg13g2_buf_2
Xfanout933 net934 net933 VPWR VGND sg13g2_buf_2
Xfanout911 net471 net911 VPWR VGND sg13g2_buf_8
Xhold497 mac1.sum_lvl2_ff\[10\] VPWR VGND net537 sg13g2_dlygate4sd3_1
Xfanout977 net281 net977 VPWR VGND sg13g2_buf_8
Xfanout944 net945 net944 VPWR VGND sg13g2_buf_8
Xfanout966 net967 net966 VPWR VGND sg13g2_buf_8
Xfanout955 DP_1.matrix\[74\] net955 VPWR VGND sg13g2_buf_8
Xfanout999 net352 net999 VPWR VGND sg13g2_buf_2
Xfanout988 net509 net988 VPWR VGND sg13g2_buf_8
X_6149_ net1059 VGND VPWR _0254_ DP_4.matrix\[38\] clknet_leaf_41_clk sg13g2_dfrbpq_1
XFILLER_9_239 VPWR VGND sg13g2_fill_1
XFILLER_10_964 VPWR VGND sg13g2_decap_8
XFILLER_6_968 VPWR VGND sg13g2_decap_8
XFILLER_49_600 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_44_393 VPWR VGND sg13g2_fill_1
X_3850_ net920 net967 net922 _0697_ VPWR VGND net965 sg13g2_nand4_1
X_3781_ _0631_ _0630_ _0623_ VPWR VGND sg13g2_nand2b_1
X_5520_ net488 _2256_ _0057_ VPWR VGND sg13g2_xor2_1
X_5451_ mac2.sum_lvl2_ff\[23\] mac2.sum_lvl2_ff\[4\] _2205_ VPWR VGND sg13g2_and2_1
X_5382_ net354 _2149_ _0026_ VPWR VGND sg13g2_xor2_1
X_4402_ _1228_ _1216_ _1229_ VPWR VGND sg13g2_xor2_1
X_4333_ _1160_ _1161_ _1162_ VPWR VGND sg13g2_and2_1
X_4264_ _1094_ _1090_ _1093_ VPWR VGND sg13g2_xnor2_1
X_3215_ _2806_ _2790_ _2804_ VPWR VGND sg13g2_xnor2_1
X_6003_ net1082 VGND VPWR _0108_ mac1.products_ff\[12\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_4195_ _1027_ _1026_ _1023_ VPWR VGND sg13g2_nand2b_1
X_3146_ _2738_ _2737_ _2734_ VPWR VGND sg13g2_nand2b_1
X_3077_ _2670_ _2637_ _2671_ VPWR VGND sg13g2_xor2_1
XFILLER_39_187 VPWR VGND sg13g2_fill_1
XFILLER_39_1000 VPWR VGND sg13g2_decap_8
XFILLER_10_216 VPWR VGND sg13g2_fill_1
XFILLER_10_238 VPWR VGND sg13g2_fill_2
X_3979_ _0823_ _0817_ _0821_ VPWR VGND sg13g2_xnor2_1
X_5718_ net771 VPWR _2426_ VGND net916 net773 sg13g2_o21ai_1
X_5649_ mac2.total_sum\[0\] mac1.total_sum\[0\] net25 VPWR VGND sg13g2_xor2_1
XFILLER_46_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_949 VPWR VGND sg13g2_decap_8
Xhold261 DP_2.matrix\[75\] VPWR VGND net301 sg13g2_dlygate4sd3_1
Xhold250 _0090_ VPWR VGND net290 sg13g2_dlygate4sd3_1
Xhold294 _0007_ VPWR VGND net334 sg13g2_dlygate4sd3_1
Xhold283 mac1.sum_lvl3_ff\[12\] VPWR VGND net323 sg13g2_dlygate4sd3_1
Xhold272 _2293_ VPWR VGND net312 sg13g2_dlygate4sd3_1
Xfanout785 net786 net785 VPWR VGND sg13g2_buf_8
Xfanout774 _2369_ net774 VPWR VGND sg13g2_buf_8
Xfanout763 _2370_ net763 VPWR VGND sg13g2_buf_8
Xfanout796 net288 net796 VPWR VGND sg13g2_buf_8
XFILLER_45_124 VPWR VGND sg13g2_fill_1
XFILLER_18_338 VPWR VGND sg13g2_fill_1
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_42_875 VPWR VGND sg13g2_decap_8
XFILLER_14_544 VPWR VGND sg13g2_decap_4
XFILLER_2_971 VPWR VGND sg13g2_decap_8
XFILLER_7_1020 VPWR VGND sg13g2_decap_8
X_3000_ _2598_ net954 net903 net898 net956 VPWR VGND sg13g2_a22oi_1
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_37_614 VPWR VGND sg13g2_decap_4
XFILLER_18_850 VPWR VGND sg13g2_fill_2
XFILLER_37_669 VPWR VGND sg13g2_fill_1
X_4951_ _1751_ _1741_ _1752_ VPWR VGND sg13g2_xor2_1
X_4882_ _1661_ _1687_ _1689_ VPWR VGND sg13g2_and2_1
X_3902_ _0748_ _0745_ _0747_ VPWR VGND sg13g2_nand2_1
X_3833_ _0681_ _0680_ _0679_ VPWR VGND sg13g2_nand2b_1
X_3764_ _0614_ _0615_ _0075_ VPWR VGND sg13g2_nor2_1
X_5503_ _0037_ _2243_ _2246_ VPWR VGND sg13g2_xnor2_1
X_6483_ net1018 VGND VPWR net426 mac2.total_sum\[11\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3695_ VGND VPWR _0552_ _0551_ _0540_ sg13g2_or2_1
X_5434_ _2193_ net409 mac1.sum_lvl3_ff\[15\] VPWR VGND sg13g2_xnor2_1
X_5365_ net265 mac1.sum_lvl2_ff\[19\] _0000_ VPWR VGND sg13g2_xor2_1
X_5296_ _2085_ mac1.sum_lvl2_ff\[20\] net332 VPWR VGND sg13g2_nand2_1
X_4316_ _1145_ _1138_ _1143_ _1144_ VPWR VGND sg13g2_and3_1
X_4247_ _1078_ _1049_ _1077_ VPWR VGND sg13g2_nand2b_1
X_4178_ _1011_ net863 net818 net865 net816 VPWR VGND sg13g2_a22oi_1
X_3129_ VGND VPWR _2718_ _2719_ _2722_ _2702_ sg13g2_a21oi_1
XFILLER_42_116 VPWR VGND sg13g2_fill_2
XFILLER_42_127 VPWR VGND sg13g2_fill_1
XFILLER_13_1003 VPWR VGND sg13g2_decap_8
XFILLER_47_967 VPWR VGND sg13g2_decap_8
XFILLER_19_658 VPWR VGND sg13g2_fill_1
XFILLER_15_897 VPWR VGND sg13g2_fill_1
XFILLER_30_878 VPWR VGND sg13g2_decap_8
X_3480_ _0343_ _0314_ _0342_ VPWR VGND sg13g2_nand2b_1
XFILLER_44_4 VPWR VGND sg13g2_fill_1
XFILLER_29_1021 VPWR VGND sg13g2_decap_8
X_5150_ _1945_ net850 net994 VPWR VGND sg13g2_nand2_1
X_5081_ _1878_ net998 net797 net839 net794 VPWR VGND sg13g2_a22oi_1
X_4101_ _0904_ _0940_ _0941_ VPWR VGND sg13g2_nor2b_1
X_4032_ _0860_ VPWR _0874_ VGND _0849_ _0861_ sg13g2_o21ai_1
XFILLER_37_411 VPWR VGND sg13g2_fill_2
XFILLER_38_956 VPWR VGND sg13g2_decap_8
XFILLER_37_455 VPWR VGND sg13g2_fill_2
X_5983_ net786 _0265_ VPWR VGND sg13g2_buf_1
XFILLER_25_639 VPWR VGND sg13g2_decap_8
XFILLER_37_488 VPWR VGND sg13g2_fill_2
X_4934_ _1736_ _1724_ _1734_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_1025 VPWR VGND sg13g2_decap_4
X_4865_ _1672_ _1643_ _1673_ VPWR VGND sg13g2_xor2_1
XFILLER_32_193 VPWR VGND sg13g2_fill_2
X_3816_ net923 net921 net969 DP_1.matrix\[41\] _0664_ VPWR VGND sg13g2_and4_1
X_4796_ _1606_ _1603_ _0139_ VPWR VGND sg13g2_xor2_1
XFILLER_20_399 VPWR VGND sg13g2_fill_2
X_3747_ _0600_ _0590_ _0602_ VPWR VGND sg13g2_xor2_1
X_3678_ _0107_ _0534_ _0535_ VPWR VGND sg13g2_xnor2_1
X_6466_ net1035 VGND VPWR _0033_ mac2.sum_lvl3_ff\[10\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5417_ _2172_ _2175_ _2179_ VPWR VGND sg13g2_nor2_1
X_6397_ net1090 VGND VPWR net184 mac2.sum_lvl1_ff\[10\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_5348_ _2124_ _2125_ _2126_ VPWR VGND sg13g2_nor2_1
XFILLER_43_1018 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
X_5279_ _2070_ _2047_ _2069_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_923 VPWR VGND sg13g2_decap_8
XFILLER_43_436 VPWR VGND sg13g2_fill_2
XFILLER_7_326 VPWR VGND sg13g2_fill_2
XFILLER_11_71 VPWR VGND sg13g2_fill_1
XFILLER_38_208 VPWR VGND sg13g2_fill_2
XFILLER_47_731 VPWR VGND sg13g2_fill_2
XFILLER_35_915 VPWR VGND sg13g2_decap_8
X_4650_ net835 net831 net874 net873 _1464_ VPWR VGND sg13g2_and4_1
X_3601_ _0460_ _0442_ _0461_ VPWR VGND sg13g2_xor2_1
Xinput10 uio_in[1] net10 VPWR VGND sg13g2_buf_1
X_6320_ net1034 VGND VPWR net48 mac2.sum_lvl3_ff\[33\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_4581_ _1397_ net827 net881 VPWR VGND sg13g2_nand2_1
X_3532_ _0393_ _0386_ _0392_ VPWR VGND sg13g2_nand2_1
X_3463_ _0297_ VPWR _0326_ VGND _0295_ _0298_ sg13g2_o21ai_1
X_6251_ net1015 VGND VPWR net43 mac1.sum_lvl1_ff\[80\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5202_ _1996_ _1986_ _1995_ VPWR VGND sg13g2_xnor2_1
X_6182_ net1067 VGND VPWR net187 mac1.sum_lvl2_ff\[3\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3394_ _2971_ _2972_ _2974_ _2975_ VPWR VGND sg13g2_nor3_1
XFILLER_35_0 VPWR VGND sg13g2_fill_1
X_5133_ _1929_ _1913_ _1928_ VPWR VGND sg13g2_nand2_1
X_5064_ _1861_ _1860_ _1857_ VPWR VGND sg13g2_nand2b_1
X_4015_ _0856_ _0857_ _0858_ VPWR VGND sg13g2_nor2b_1
X_5966_ net271 _0240_ VPWR VGND sg13g2_buf_1
XFILLER_12_108 VPWR VGND sg13g2_fill_1
X_4917_ _1720_ net851 net799 net796 net853 VPWR VGND sg13g2_a22oi_1
X_5897_ _2576_ net827 net759 VPWR VGND sg13g2_nand2_1
X_4848_ _1654_ _1653_ _1657_ VPWR VGND sg13g2_xor2_1
XFILLER_21_664 VPWR VGND sg13g2_fill_1
X_4779_ _1586_ _1588_ _1589_ _1590_ VPWR VGND sg13g2_nor3_1
XFILLER_5_819 VPWR VGND sg13g2_decap_4
XFILLER_10_1006 VPWR VGND sg13g2_decap_8
X_6449_ net1090 VGND VPWR net125 mac2.sum_lvl2_ff\[28\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_44_789 VPWR VGND sg13g2_fill_1
XFILLER_40_962 VPWR VGND sg13g2_decap_8
XFILLER_7_167 VPWR VGND sg13g2_fill_2
XFILLER_4_896 VPWR VGND sg13g2_fill_2
XFILLER_26_1013 VPWR VGND sg13g2_decap_8
XFILLER_19_285 VPWR VGND sg13g2_fill_1
X_5820_ VGND VPWR net996 net760 _2526_ _2525_ sg13g2_a21oi_1
XFILLER_16_970 VPWR VGND sg13g2_decap_8
X_5751_ _2455_ VPWR _2458_ VGND _2456_ _2457_ sg13g2_o21ai_1
XFILLER_31_962 VPWR VGND sg13g2_decap_8
X_4702_ _1504_ _1512_ _1514_ _1515_ VPWR VGND sg13g2_or3_1
X_5682_ net770 VPWR _2391_ VGND net973 net773 sg13g2_o21ai_1
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_61 VPWR VGND sg13g2_fill_1
X_4633_ _1447_ _1446_ _0145_ VPWR VGND sg13g2_xor2_1
X_4564_ _1379_ _1380_ _1374_ _1381_ VPWR VGND sg13g2_nand3_1
X_3515_ _0353_ VPWR _0377_ VGND _0373_ _0375_ sg13g2_o21ai_1
X_6303_ net1024 VGND VPWR _0003_ mac1.sum_lvl3_ff\[12\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_4495_ _1316_ _1299_ _1319_ VPWR VGND sg13g2_xor2_1
X_6234_ net1035 VGND VPWR net222 mac2.sum_lvl2_ff\[45\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3446_ _0306_ _0307_ _0270_ _0310_ VPWR VGND sg13g2_nand3_1
X_3377_ net993 net937 _0069_ VPWR VGND sg13g2_and2_1
X_6165_ net1064 VGND VPWR net231 mac1.sum_lvl1_ff\[38\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_6096_ net1046 VGND VPWR _0217_ DP_2.matrix\[77\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5116_ _1910_ _1902_ _1912_ VPWR VGND sg13g2_xor2_1
X_5047_ VGND VPWR _1841_ _1842_ _1845_ _1824_ sg13g2_a21oi_1
XFILLER_38_550 VPWR VGND sg13g2_fill_1
X_5949_ net895 _0215_ VPWR VGND sg13g2_buf_1
XFILLER_40_203 VPWR VGND sg13g2_fill_1
XFILLER_41_759 VPWR VGND sg13g2_fill_2
XFILLER_22_962 VPWR VGND sg13g2_decap_8
XFILLER_49_1024 VPWR VGND sg13g2_decap_4
XFILLER_1_899 VPWR VGND sg13g2_decap_8
XFILLER_1_1004 VPWR VGND sg13g2_decap_8
XFILLER_29_594 VPWR VGND sg13g2_fill_2
XFILLER_32_704 VPWR VGND sg13g2_fill_1
XFILLER_32_748 VPWR VGND sg13g2_fill_1
XFILLER_8_443 VPWR VGND sg13g2_fill_1
XFILLER_9_966 VPWR VGND sg13g2_decap_8
X_3300_ _2858_ VPWR _2888_ VGND _2856_ _2859_ sg13g2_o21ai_1
X_4280_ _1088_ _1107_ _1109_ _1110_ VPWR VGND sg13g2_or3_1
X_3231_ _2821_ net955 net1003 VPWR VGND sg13g2_nand2_1
X_3162_ net900 net941 net905 _2754_ VPWR VGND net1006 sg13g2_nand4_1
XFILLER_12_2 VPWR VGND sg13g2_fill_1
XFILLER_48_870 VPWR VGND sg13g2_decap_8
X_3093_ VGND VPWR _2684_ _2685_ _2687_ _2667_ sg13g2_a21oi_1
X_5803_ _2508_ _2506_ _2509_ VPWR VGND sg13g2_nor2b_1
X_3995_ _0825_ VPWR _0838_ VGND _0809_ _0826_ sg13g2_o21ai_1
X_5734_ _2591_ _2411_ net755 _2442_ VPWR VGND sg13g2_mux2_1
X_5665_ VGND VPWR _2590_ net773 _2374_ _2373_ sg13g2_a21oi_1
X_4616_ net831 net876 net836 _1431_ VPWR VGND net874 sg13g2_nand4_1
X_5596_ VGND VPWR _2314_ _2316_ _2317_ _2315_ sg13g2_a21oi_1
Xhold410 _0043_ VPWR VGND net450 sg13g2_dlygate4sd3_1
Xhold432 DP_3.matrix\[42\] VPWR VGND net472 sg13g2_dlygate4sd3_1
Xhold443 mac1.sum_lvl3_ff\[6\] VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold454 mac1.sum_lvl2_ff\[3\] VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold421 mac2.sum_lvl2_ff\[4\] VPWR VGND net461 sg13g2_dlygate4sd3_1
X_4547_ _1365_ _1364_ _1357_ VPWR VGND sg13g2_nand2b_1
X_4478_ _1302_ net861 net995 VPWR VGND sg13g2_nand2_1
Xhold476 _2104_ VPWR VGND net516 sg13g2_dlygate4sd3_1
Xhold465 DP_1.matrix\[7\] VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold487 _0044_ VPWR VGND net527 sg13g2_dlygate4sd3_1
X_3429_ _0291_ _0288_ _0293_ VPWR VGND sg13g2_xor2_1
X_6217_ net1022 VGND VPWR net201 mac1.sum_lvl2_ff\[44\] clknet_leaf_0_clk sg13g2_dfrbpq_1
Xfanout901 net902 net901 VPWR VGND sg13g2_buf_1
Xfanout923 net391 net923 VPWR VGND sg13g2_buf_2
Xfanout934 net935 net934 VPWR VGND sg13g2_buf_1
Xfanout912 net913 net912 VPWR VGND sg13g2_buf_8
Xhold498 _2116_ VPWR VGND net538 sg13g2_dlygate4sd3_1
Xfanout956 net957 net956 VPWR VGND sg13g2_buf_8
Xfanout967 net522 net967 VPWR VGND sg13g2_buf_8
Xfanout945 DP_1.matrix\[78\] net945 VPWR VGND sg13g2_buf_8
X_6148_ net1060 VGND VPWR _0253_ DP_4.matrix\[37\] clknet_leaf_31_clk sg13g2_dfrbpq_2
Xfanout989 net402 net989 VPWR VGND sg13g2_buf_8
Xfanout978 net979 net978 VPWR VGND sg13g2_buf_2
X_6079_ net1019 VGND VPWR _0095_ mac1.products_ff\[146\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_39_881 VPWR VGND sg13g2_decap_8
XFILLER_9_218 VPWR VGND sg13g2_fill_2
XFILLER_13_269 VPWR VGND sg13g2_fill_2
XFILLER_16_1012 VPWR VGND sg13g2_decap_8
XFILLER_10_943 VPWR VGND sg13g2_decap_8
XFILLER_6_947 VPWR VGND sg13g2_decap_8
XFILLER_23_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_656 VPWR VGND sg13g2_decap_4
XFILLER_37_807 VPWR VGND sg13g2_fill_1
XFILLER_17_564 VPWR VGND sg13g2_fill_1
XFILLER_45_895 VPWR VGND sg13g2_decap_8
X_3780_ _0628_ _0629_ _0630_ VPWR VGND sg13g2_nor2b_1
XFILLER_12_291 VPWR VGND sg13g2_fill_1
X_5450_ _2202_ VPWR _2204_ VGND _2201_ _2203_ sg13g2_o21ai_1
X_4401_ _1226_ _1217_ _1228_ VPWR VGND sg13g2_xor2_1
X_5381_ net353 mac1.sum_lvl3_ff\[24\] _2151_ VPWR VGND sg13g2_xor2_1
X_4332_ _1158_ _1157_ _1159_ _1161_ VPWR VGND sg13g2_a21o_1
X_4263_ _1093_ _1056_ _1091_ VPWR VGND sg13g2_xnor2_1
X_3214_ _2805_ _2790_ _2804_ VPWR VGND sg13g2_nand2_1
X_6002_ net1070 VGND VPWR _0107_ mac1.products_ff\[11\] clknet_leaf_44_clk sg13g2_dfrbpq_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
X_4194_ _1025_ _1004_ _1026_ VPWR VGND sg13g2_xor2_1
X_3145_ _2736_ _2697_ _2737_ VPWR VGND sg13g2_xor2_1
X_3076_ _2670_ net952 net894 VPWR VGND sg13g2_nand2_1
XFILLER_35_383 VPWR VGND sg13g2_fill_2
X_3978_ _0822_ _0817_ _0821_ VPWR VGND sg13g2_nand2_1
X_5717_ _2425_ net897 net763 VPWR VGND sg13g2_nand2_1
X_5648_ net24 _2357_ _2358_ VPWR VGND sg13g2_xnor2_1
X_5579_ _2304_ mac1.total_sum\[0\] mac2.total_sum\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_3_928 VPWR VGND sg13g2_decap_8
Xhold240 DP_2.matrix\[78\] VPWR VGND net280 sg13g2_dlygate4sd3_1
Xhold251 mac2.sum_lvl2_ff\[19\] VPWR VGND net291 sg13g2_dlygate4sd3_1
Xhold262 DP_3.matrix\[74\] VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold295 DP_2.matrix\[38\] VPWR VGND net335 sg13g2_dlygate4sd3_1
Xhold284 _2183_ VPWR VGND net324 sg13g2_dlygate4sd3_1
Xhold273 _0051_ VPWR VGND net313 sg13g2_dlygate4sd3_1
Xfanout753 net754 net753 VPWR VGND sg13g2_buf_8
Xfanout775 net776 net775 VPWR VGND sg13g2_buf_8
Xfanout764 _2370_ net764 VPWR VGND sg13g2_buf_8
Xfanout786 net356 net786 VPWR VGND sg13g2_buf_1
Xfanout797 net798 net797 VPWR VGND sg13g2_buf_2
XFILLER_19_829 VPWR VGND sg13g2_fill_2
XFILLER_46_648 VPWR VGND sg13g2_fill_2
XFILLER_41_331 VPWR VGND sg13g2_fill_1
XFILLER_6_777 VPWR VGND sg13g2_fill_2
XFILLER_2_950 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_17_350 VPWR VGND sg13g2_decap_8
X_4950_ _1751_ _1749_ _1750_ VPWR VGND sg13g2_nand2_1
X_4881_ _1688_ _1687_ _0142_ VPWR VGND sg13g2_xor2_1
X_3901_ _0744_ _0743_ _0714_ _0747_ VPWR VGND sg13g2_a21o_1
X_3832_ _0652_ VPWR _0680_ VGND _0676_ _0677_ sg13g2_o21ai_1
XFILLER_20_526 VPWR VGND sg13g2_fill_1
X_5502_ mac2.sum_lvl2_ff\[14\] mac2.sum_lvl2_ff\[33\] _2246_ VPWR VGND sg13g2_xor2_1
X_3763_ _0615_ net918 net977 net975 net924 VPWR VGND sg13g2_a22oi_1
X_6482_ net1017 VGND VPWR net382 mac2.total_sum\[10\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3694_ _0549_ _0541_ _0551_ VPWR VGND sg13g2_xor2_1
X_5433_ _2188_ VPWR _2192_ VGND _2189_ _2191_ sg13g2_o21ai_1
XFILLER_10_29 VPWR VGND sg13g2_fill_1
X_5364_ _0006_ _2137_ net286 VPWR VGND sg13g2_xnor2_1
X_4315_ _1139_ VPWR _1144_ VGND _1140_ _1142_ sg13g2_o21ai_1
X_5295_ _2084_ mac1.sum_lvl2_ff\[19\] net265 VPWR VGND sg13g2_nand2_1
X_4246_ _1077_ _1053_ _1076_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_604 VPWR VGND sg13g2_fill_1
X_4177_ net816 net865 net818 _1010_ VPWR VGND net863 sg13g2_nand4_1
X_3128_ _2718_ _2719_ _2702_ _2721_ VPWR VGND sg13g2_nand3_1
X_3059_ _2652_ _2653_ _2635_ _2654_ VPWR VGND sg13g2_nand3_1
XFILLER_36_681 VPWR VGND sg13g2_fill_2
XFILLER_23_364 VPWR VGND sg13g2_fill_2
XFILLER_24_887 VPWR VGND sg13g2_fill_1
XFILLER_3_758 VPWR VGND sg13g2_fill_1
XFILLER_47_946 VPWR VGND sg13g2_decap_8
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_29_1000 VPWR VGND sg13g2_decap_8
X_5080_ net793 net839 net798 _1877_ VPWR VGND net998 sg13g2_nand4_1
X_4100_ _0940_ _0935_ _0938_ VPWR VGND sg13g2_xnor2_1
X_4031_ _0846_ _0840_ _0848_ _0873_ VPWR VGND sg13g2_a21o_1
XFILLER_38_935 VPWR VGND sg13g2_decap_8
X_5982_ net788 _0264_ VPWR VGND sg13g2_buf_1
X_4933_ _1735_ _1734_ _1724_ VPWR VGND sg13g2_nand2b_1
XFILLER_33_662 VPWR VGND sg13g2_fill_2
XFILLER_33_673 VPWR VGND sg13g2_fill_2
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
X_4864_ _1672_ net821 DP_3.matrix\[7\] VPWR VGND sg13g2_nand2_1
X_3815_ _0663_ net917 net971 VPWR VGND sg13g2_nand2_1
X_4795_ _1606_ _1604_ _1605_ VPWR VGND sg13g2_nand2b_1
X_3746_ _0600_ _0590_ _0601_ VPWR VGND sg13g2_nor2b_1
X_6465_ net1035 VGND VPWR _0047_ mac2.sum_lvl3_ff\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5416_ _2173_ _2176_ _2178_ VPWR VGND sg13g2_nor2_1
X_3677_ VGND VPWR _0502_ _0505_ _0535_ _0500_ sg13g2_a21oi_1
X_6396_ net1089 VGND VPWR net228 mac2.sum_lvl1_ff\[9\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5347_ _2120_ _2115_ _2119_ _2125_ VPWR VGND sg13g2_a21o_1
X_5278_ _2067_ _2066_ _2069_ VPWR VGND sg13g2_xor2_1
XFILLER_29_902 VPWR VGND sg13g2_decap_8
X_4229_ _1060_ _1055_ _1058_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_979 VPWR VGND sg13g2_decap_8
XFILLER_44_949 VPWR VGND sg13g2_decap_8
XFILLER_8_806 VPWR VGND sg13g2_fill_2
XFILLER_7_305 VPWR VGND sg13g2_fill_1
XFILLER_12_879 VPWR VGND sg13g2_fill_1
XFILLER_20_890 VPWR VGND sg13g2_fill_2
XFILLER_3_522 VPWR VGND sg13g2_fill_2
XFILLER_47_721 VPWR VGND sg13g2_fill_1
XFILLER_4_1024 VPWR VGND sg13g2_decap_4
XFILLER_47_765 VPWR VGND sg13g2_decap_8
XFILLER_47_776 VPWR VGND sg13g2_fill_1
XFILLER_34_448 VPWR VGND sg13g2_fill_2
XFILLER_15_673 VPWR VGND sg13g2_fill_1
X_3600_ _0460_ _0443_ _0458_ VPWR VGND sg13g2_xnor2_1
X_4580_ _1377_ VPWR _1396_ VGND _1375_ _1378_ sg13g2_o21ai_1
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
X_3531_ _0392_ _0387_ _0390_ VPWR VGND sg13g2_xnor2_1
X_6250_ net1015 VGND VPWR net166 mac1.sum_lvl1_ff\[79\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3462_ _0325_ _0320_ _0323_ VPWR VGND sg13g2_xnor2_1
X_5201_ _1995_ _1987_ _1993_ VPWR VGND sg13g2_xnor2_1
X_3393_ _2974_ net987 net937 net989 net932 VPWR VGND sg13g2_a22oi_1
X_6181_ net1064 VGND VPWR net114 mac1.sum_lvl2_ff\[2\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_5132_ _1927_ _1920_ _1928_ VPWR VGND sg13g2_xor2_1
X_5063_ _1859_ _1819_ _1860_ VPWR VGND sg13g2_xor2_1
X_4014_ _0852_ VPWR _0857_ VGND _0854_ _0855_ sg13g2_o21ai_1
XFILLER_38_776 VPWR VGND sg13g2_decap_8
X_5965_ net849 _0239_ VPWR VGND sg13g2_buf_1
XFILLER_33_481 VPWR VGND sg13g2_fill_1
XFILLER_34_982 VPWR VGND sg13g2_decap_8
X_4916_ net799 net853 net796 net851 _1719_ VPWR VGND sg13g2_and4_1
X_5896_ _2508_ _2506_ _2575_ VPWR VGND sg13g2_xor2_1
X_4847_ _1653_ _1654_ _1656_ VPWR VGND sg13g2_nor2b_1
X_4778_ _1589_ net872 net826 net875 net823 VPWR VGND sg13g2_a22oi_1
X_3729_ _0585_ _0565_ _0582_ VPWR VGND sg13g2_xnor2_1
X_6448_ net1089 VGND VPWR net88 mac2.sum_lvl2_ff\[27\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6379_ net1027 VGND VPWR _0158_ mac2.products_ff\[144\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_44_746 VPWR VGND sg13g2_fill_2
XFILLER_8_603 VPWR VGND sg13g2_fill_2
XFILLER_24_492 VPWR VGND sg13g2_fill_1
XFILLER_40_941 VPWR VGND sg13g2_decap_8
XFILLER_22_82 VPWR VGND sg13g2_fill_1
XFILLER_47_562 VPWR VGND sg13g2_decap_4
X_5750_ net768 VPWR _2457_ VGND net876 net777 sg13g2_o21ai_1
XFILLER_22_418 VPWR VGND sg13g2_fill_2
X_5681_ _2390_ net276 net763 VPWR VGND sg13g2_nand2_1
XFILLER_31_941 VPWR VGND sg13g2_decap_8
XFILLER_33_1007 VPWR VGND sg13g2_decap_8
X_4701_ VGND VPWR _1510_ _1511_ _1514_ _1505_ sg13g2_a21oi_1
X_4632_ VGND VPWR _1388_ _1414_ _1447_ _1413_ sg13g2_a21oi_1
X_4563_ _1375_ VPWR _1380_ VGND _1376_ _1378_ sg13g2_o21ai_1
X_4494_ _1299_ _1316_ _1318_ VPWR VGND sg13g2_nor2_1
X_3514_ _0353_ _0373_ _0375_ _0376_ VPWR VGND sg13g2_or3_1
X_6302_ net1024 VGND VPWR _0002_ mac1.sum_lvl3_ff\[11\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_3445_ _0309_ _0270_ _0306_ _0307_ VPWR VGND sg13g2_and3_1
X_6233_ net1036 VGND VPWR net190 mac2.sum_lvl2_ff\[44\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6164_ net1045 VGND VPWR net92 mac1.sum_lvl1_ff\[37\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3376_ _0100_ _2953_ _2960_ VPWR VGND sg13g2_xnor2_1
X_6095_ net1042 VGND VPWR _0216_ DP_2.matrix\[76\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5115_ _1910_ _1902_ _1911_ VPWR VGND sg13g2_nor2b_1
X_5046_ _1841_ _1842_ _1824_ _1844_ VPWR VGND sg13g2_nand3_1
XFILLER_25_201 VPWR VGND sg13g2_fill_1
XFILLER_26_746 VPWR VGND sg13g2_fill_1
XFILLER_41_716 VPWR VGND sg13g2_fill_1
X_5948_ net897 _0214_ VPWR VGND sg13g2_buf_1
XFILLER_13_429 VPWR VGND sg13g2_fill_2
X_5879_ _2564_ VPWR _0223_ VGND net759 _2563_ sg13g2_o21ai_1
XFILLER_49_1003 VPWR VGND sg13g2_decap_8
XFILLER_9_945 VPWR VGND sg13g2_decap_8
XFILLER_13_996 VPWR VGND sg13g2_decap_8
XFILLER_8_488 VPWR VGND sg13g2_fill_2
XFILLER_4_661 VPWR VGND sg13g2_fill_1
XFILLER_3_171 VPWR VGND sg13g2_fill_2
X_3230_ _2793_ VPWR _2820_ VGND _2791_ _2794_ sg13g2_o21ai_1
X_3161_ net905 net900 net941 net1006 _2753_ VPWR VGND sg13g2_and4_1
X_3092_ _2684_ _2685_ _2667_ _2686_ VPWR VGND sg13g2_nand3_1
X_5802_ _2508_ _2507_ net769 net765 net792 VPWR VGND sg13g2_a22oi_1
X_3994_ _0806_ _0800_ _0808_ _0837_ VPWR VGND sg13g2_a21o_1
X_5733_ _2441_ net772 _2440_ net764 net888 VPWR VGND sg13g2_a22oi_1
X_5664_ net771 VPWR _2373_ VGND DP_1.matrix\[44\] _2369_ sg13g2_o21ai_1
X_5595_ _2316_ _2314_ net29 VPWR VGND sg13g2_xor2_1
X_4615_ net835 net832 net876 net874 _1430_ VPWR VGND sg13g2_and4_1
Xhold411 mac2.sum_lvl3_ff\[2\] VPWR VGND net451 sg13g2_dlygate4sd3_1
Xhold400 DP_4.matrix\[37\] VPWR VGND net440 sg13g2_dlygate4sd3_1
X_4546_ _1362_ _1363_ _1364_ VPWR VGND sg13g2_nor2b_1
Xhold444 _2156_ VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold422 _2206_ VPWR VGND net462 sg13g2_dlygate4sd3_1
Xhold433 DP_3.matrix\[39\] VPWR VGND net473 sg13g2_dlygate4sd3_1
X_4477_ _1280_ VPWR _1301_ VGND _1252_ _1278_ sg13g2_o21ai_1
Xhold477 DP_3.matrix\[4\] VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold455 _2093_ VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold466 mac2.sum_lvl2_ff\[7\] VPWR VGND net506 sg13g2_dlygate4sd3_1
X_3428_ _0292_ _0291_ _0288_ VPWR VGND sg13g2_nand2b_1
Xfanout902 net345 net902 VPWR VGND sg13g2_buf_1
Xfanout924 net391 net924 VPWR VGND sg13g2_buf_8
X_6216_ net1022 VGND VPWR net153 mac1.sum_lvl2_ff\[43\] clknet_leaf_66_clk sg13g2_dfrbpq_1
Xfanout913 net523 net913 VPWR VGND sg13g2_buf_8
Xhold488 DP_1.matrix\[42\] VPWR VGND net528 sg13g2_dlygate4sd3_1
Xhold499 mac2.sum_lvl3_ff\[7\] VPWR VGND net539 sg13g2_dlygate4sd3_1
Xfanout935 net936 net935 VPWR VGND sg13g2_buf_1
Xfanout946 net947 net946 VPWR VGND sg13g2_buf_2
Xfanout968 net969 net968 VPWR VGND sg13g2_buf_8
Xfanout957 net304 net957 VPWR VGND sg13g2_buf_8
X_3359_ _2919_ VPWR _2945_ VGND _2890_ _2917_ sg13g2_o21ai_1
X_6147_ net1060 VGND VPWR _0252_ DP_4.matrix\[36\] clknet_leaf_31_clk sg13g2_dfrbpq_2
Xfanout979 net980 net979 VPWR VGND sg13g2_buf_1
X_6078_ net1086 VGND VPWR _0205_ DP_2.matrix\[37\] clknet_leaf_50_clk sg13g2_dfrbpq_2
XFILLER_39_860 VPWR VGND sg13g2_decap_8
X_5029_ _1827_ net789 net846 VPWR VGND sg13g2_nand2_1
XFILLER_41_557 VPWR VGND sg13g2_decap_4
XFILLER_6_926 VPWR VGND sg13g2_decap_8
XFILLER_10_999 VPWR VGND sg13g2_decap_8
XFILLER_49_635 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_45_874 VPWR VGND sg13g2_decap_8
XFILLER_17_587 VPWR VGND sg13g2_fill_1
XFILLER_12_270 VPWR VGND sg13g2_fill_2
X_4400_ _1227_ _1217_ _1226_ VPWR VGND sg13g2_nand2b_1
X_5380_ mac1.sum_lvl3_ff\[24\] mac1.sum_lvl3_ff\[4\] _2150_ VPWR VGND sg13g2_and2_1
XFILLER_5_63 VPWR VGND sg13g2_fill_1
X_4331_ _1158_ _1159_ _1157_ _1160_ VPWR VGND sg13g2_nand3_1
X_4262_ VGND VPWR _1092_ _1091_ _1056_ sg13g2_or2_1
X_3213_ _2803_ _2796_ _2804_ VPWR VGND sg13g2_xor2_1
X_6001_ net1070 VGND VPWR _0106_ mac1.products_ff\[10\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_4193_ _1025_ net868 net809 VPWR VGND sg13g2_nand2_1
X_3144_ _2736_ net955 net889 VPWR VGND sg13g2_nand2_1
X_3075_ _2669_ net953 net892 VPWR VGND sg13g2_nand2_1
XFILLER_35_373 VPWR VGND sg13g2_fill_1
XFILLER_36_885 VPWR VGND sg13g2_decap_8
X_3977_ _0819_ _0820_ _0821_ VPWR VGND sg13g2_nor2_1
XFILLER_23_579 VPWR VGND sg13g2_fill_2
X_5716_ _2424_ _2423_ _2419_ VPWR VGND sg13g2_nand2b_1
X_5647_ _2358_ mac1.total_sum\[15\] mac2.total_sum\[15\] VPWR VGND sg13g2_xnor2_1
XFILLER_40_38 VPWR VGND sg13g2_decap_8
X_5578_ net305 mac2.sum_lvl3_ff\[20\] _0048_ VPWR VGND sg13g2_xor2_1
Xhold241 DP_1.matrix\[36\] VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold230 DP_1.matrix\[79\] VPWR VGND net270 sg13g2_dlygate4sd3_1
Xhold252 _0039_ VPWR VGND net292 sg13g2_dlygate4sd3_1
X_4529_ _1349_ net829 net886 net884 net833 VPWR VGND sg13g2_a22oi_1
Xhold263 DP_4.matrix\[74\] VPWR VGND net303 sg13g2_dlygate4sd3_1
Xhold296 DP_1.matrix\[77\] VPWR VGND net336 sg13g2_dlygate4sd3_1
Xhold285 _0019_ VPWR VGND net325 sg13g2_dlygate4sd3_1
Xhold274 DP_4.matrix\[40\] VPWR VGND net314 sg13g2_dlygate4sd3_1
Xfanout765 net766 net765 VPWR VGND sg13g2_buf_8
Xfanout754 net757 net754 VPWR VGND sg13g2_buf_8
Xfanout776 _2368_ net776 VPWR VGND sg13g2_buf_8
Xfanout798 net800 net798 VPWR VGND sg13g2_buf_1
Xfanout787 net788 net787 VPWR VGND sg13g2_buf_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_14_557 VPWR VGND sg13g2_fill_1
Xinput9 uio_in[0] net9 VPWR VGND sg13g2_buf_1
XFILLER_18_852 VPWR VGND sg13g2_fill_1
X_4880_ _1688_ _1660_ _1666_ VPWR VGND sg13g2_nand2_1
XFILLER_44_170 VPWR VGND sg13g2_fill_1
X_3900_ VGND VPWR _0743_ _0744_ _0746_ _0714_ sg13g2_a21oi_1
XFILLER_32_310 VPWR VGND sg13g2_fill_1
XFILLER_33_855 VPWR VGND sg13g2_fill_2
X_3831_ _0652_ _0676_ _0677_ _0679_ VPWR VGND sg13g2_nor3_1
XFILLER_32_343 VPWR VGND sg13g2_fill_2
XFILLER_33_888 VPWR VGND sg13g2_decap_8
X_3762_ _0614_ net975 net918 _0074_ VPWR VGND sg13g2_and3_2
X_5501_ mac2.sum_lvl2_ff\[33\] mac2.sum_lvl2_ff\[14\] _2245_ VPWR VGND sg13g2_nor2_1
X_3693_ _0549_ _0541_ _0550_ VPWR VGND sg13g2_nor2b_1
X_6481_ net1017 VGND VPWR net340 mac2.total_sum\[9\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5432_ _0021_ net374 _2191_ VPWR VGND sg13g2_xnor2_1
X_5363_ _2138_ mac1.sum_lvl2_ff\[34\] net285 VPWR VGND sg13g2_xnor2_1
X_4314_ _1139_ _1140_ _1142_ _1143_ VPWR VGND sg13g2_or3_1
X_5294_ _0155_ _2076_ _2083_ VPWR VGND sg13g2_xnor2_1
X_4245_ _1076_ _1073_ _1075_ VPWR VGND sg13g2_nand2_1
X_4176_ net818 net816 net865 net863 _1009_ VPWR VGND sg13g2_and4_1
X_3127_ _2720_ _2702_ _2718_ _2719_ VPWR VGND sg13g2_and3_1
X_3058_ _2641_ VPWR _2653_ VGND _2649_ _2651_ sg13g2_o21ai_1
XFILLER_42_118 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_62_clk clknet_4_2_0_clk clknet_leaf_62_clk VPWR VGND sg13g2_buf_8
XFILLER_35_192 VPWR VGND sg13g2_fill_2
XFILLER_47_925 VPWR VGND sg13g2_decap_8
XFILLER_19_616 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_53_clk clknet_4_10_0_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
XFILLER_41_162 VPWR VGND sg13g2_fill_2
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
X_4030_ _0872_ _0869_ _0117_ VPWR VGND sg13g2_xor2_1
XFILLER_38_914 VPWR VGND sg13g2_decap_8
XFILLER_37_413 VPWR VGND sg13g2_fill_1
XFILLER_37_435 VPWR VGND sg13g2_fill_1
XFILLER_37_457 VPWR VGND sg13g2_fill_1
X_5981_ net790 _0263_ VPWR VGND sg13g2_buf_1
XFILLER_46_980 VPWR VGND sg13g2_decap_8
XFILLER_45_490 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_44_clk clknet_4_11_0_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
X_4932_ _1734_ _1725_ _1732_ VPWR VGND sg13g2_xnor2_1
X_4863_ _1671_ net872 net820 VPWR VGND sg13g2_nand2_1
XFILLER_21_836 VPWR VGND sg13g2_fill_1
X_3814_ _0643_ VPWR _0662_ VGND _0641_ _0644_ sg13g2_o21ai_1
XFILLER_21_869 VPWR VGND sg13g2_fill_1
X_4794_ VGND VPWR _1527_ _1567_ _1605_ _1568_ sg13g2_a21oi_1
X_3745_ _0600_ _0577_ _0599_ VPWR VGND sg13g2_xnor2_1
X_6464_ net1035 VGND VPWR net508 mac2.sum_lvl3_ff\[8\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5415_ _0018_ net394 _2177_ VPWR VGND sg13g2_xnor2_1
X_3676_ _0532_ _0533_ _0534_ VPWR VGND sg13g2_nor2b_1
X_6395_ net1089 VGND VPWR net111 mac2.sum_lvl1_ff\[8\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5346_ _2113_ _2117_ _2123_ _2124_ VPWR VGND sg13g2_nor3_1
X_5277_ _2068_ _2066_ _2067_ VPWR VGND sg13g2_nand2_1
X_4228_ _1059_ _1058_ _1055_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_446 VPWR VGND sg13g2_fill_1
XFILLER_29_958 VPWR VGND sg13g2_decap_8
X_4159_ net813 net867 net818 _0993_ VPWR VGND net865 sg13g2_nand4_1
XFILLER_44_928 VPWR VGND sg13g2_decap_8
XFILLER_16_619 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_35_clk clknet_4_15_0_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_7_328 VPWR VGND sg13g2_fill_1
XFILLER_11_40 VPWR VGND sg13g2_fill_2
XFILLER_4_1003 VPWR VGND sg13g2_decap_8
XFILLER_34_438 VPWR VGND sg13g2_fill_2
XFILLER_36_81 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_26_clk clknet_4_7_0_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_43_983 VPWR VGND sg13g2_decap_8
Xinput12 uio_in[3] net12 VPWR VGND sg13g2_buf_1
X_3530_ _0391_ _0390_ _0387_ VPWR VGND sg13g2_nand2b_1
X_3461_ _0324_ _0323_ _0320_ VPWR VGND sg13g2_nand2b_1
X_5200_ _1994_ _1987_ _1993_ VPWR VGND sg13g2_nand2_1
X_3392_ net932 net989 net940 _2973_ VPWR VGND net987 sg13g2_nand4_1
X_6180_ net1045 VGND VPWR net205 mac1.sum_lvl2_ff\[1\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5131_ _1927_ _1921_ _1925_ VPWR VGND sg13g2_xnor2_1
X_5062_ _1859_ net850 net783 VPWR VGND sg13g2_nand2_1
X_4013_ _0852_ _0854_ _0855_ _0856_ VPWR VGND sg13g2_nor3_1
XFILLER_19_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_4_4_0_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_34_961 VPWR VGND sg13g2_decap_8
X_5964_ net851 _0238_ VPWR VGND sg13g2_buf_1
X_5895_ _2574_ VPWR _0245_ VGND net758 _2573_ sg13g2_o21ai_1
X_4915_ net854 net792 _1718_ VPWR VGND sg13g2_and2_1
X_4846_ _1655_ _1653_ _1654_ VPWR VGND sg13g2_nand2b_1
XFILLER_20_110 VPWR VGND sg13g2_fill_1
XFILLER_20_132 VPWR VGND sg13g2_fill_2
XFILLER_21_644 VPWR VGND sg13g2_fill_1
X_4777_ net825 net823 net875 DP_3.matrix\[7\] _1588_ VPWR VGND sg13g2_and4_1
X_3728_ _0582_ _0565_ _0584_ VPWR VGND sg13g2_nor2b_1
X_3659_ _0489_ VPWR _0517_ VGND _0486_ _0490_ sg13g2_o21ai_1
X_6447_ net1081 VGND VPWR net156 mac2.sum_lvl2_ff\[26\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6378_ net1035 VGND VPWR _0157_ mac2.products_ff\[143\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5329_ _2107_ _2109_ net500 _2111_ VPWR VGND sg13g2_nand3_1
XFILLER_29_722 VPWR VGND sg13g2_fill_2
XFILLER_19_1022 VPWR VGND sg13g2_decap_8
XFILLER_25_994 VPWR VGND sg13g2_decap_8
XFILLER_40_920 VPWR VGND sg13g2_decap_8
XFILLER_8_637 VPWR VGND sg13g2_fill_2
XFILLER_12_666 VPWR VGND sg13g2_fill_2
XFILLER_40_997 VPWR VGND sg13g2_decap_8
XFILLER_11_198 VPWR VGND sg13g2_fill_1
XFILLER_7_169 VPWR VGND sg13g2_fill_1
XFILLER_3_375 VPWR VGND sg13g2_fill_2
XFILLER_35_736 VPWR VGND sg13g2_fill_2
XFILLER_31_920 VPWR VGND sg13g2_decap_8
X_5680_ _2389_ _2388_ _2384_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_493 VPWR VGND sg13g2_fill_1
X_4700_ _1510_ _1511_ _1505_ _1513_ VPWR VGND sg13g2_nand3_1
XFILLER_31_997 VPWR VGND sg13g2_decap_8
X_4631_ _1444_ _1416_ _1446_ VPWR VGND sg13g2_xor2_1
X_4562_ _1375_ _1376_ _1378_ _1379_ VPWR VGND sg13g2_or3_1
X_4493_ _1317_ _1299_ _1316_ VPWR VGND sg13g2_nand2_1
X_3513_ VGND VPWR _0371_ _0372_ _0375_ _0354_ sg13g2_a21oi_1
X_6301_ net1024 VGND VPWR _0001_ mac1.sum_lvl3_ff\[10\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3444_ VGND VPWR _0306_ _0307_ _0308_ _0270_ sg13g2_a21oi_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_6232_ net1049 VGND VPWR net194 mac2.sum_lvl2_ff\[43\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_6163_ net1043 VGND VPWR net224 mac1.sum_lvl1_ff\[36\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3375_ _2960_ _2954_ _2959_ VPWR VGND sg13g2_xnor2_1
X_6094_ net1046 VGND VPWR _0100_ mac1.products_ff\[151\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5114_ _1910_ _1903_ _1909_ VPWR VGND sg13g2_xnor2_1
X_5045_ _1843_ _1824_ _1841_ _1842_ VPWR VGND sg13g2_and3_1
XFILLER_26_703 VPWR VGND sg13g2_decap_8
XFILLER_26_714 VPWR VGND sg13g2_fill_1
XFILLER_38_563 VPWR VGND sg13g2_fill_1
X_5947_ net902 _0213_ VPWR VGND sg13g2_buf_1
XFILLER_22_997 VPWR VGND sg13g2_decap_8
X_5878_ _2564_ net880 net759 VPWR VGND sg13g2_nand2_1
X_4829_ VGND VPWR _1638_ _1637_ _1587_ sg13g2_or2_1
XFILLER_21_474 VPWR VGND sg13g2_fill_1
XFILLER_5_618 VPWR VGND sg13g2_fill_1
XFILLER_0_367 VPWR VGND sg13g2_fill_1
XFILLER_29_596 VPWR VGND sg13g2_fill_1
XFILLER_44_544 VPWR VGND sg13g2_fill_1
XFILLER_13_975 VPWR VGND sg13g2_decap_8
XFILLER_40_794 VPWR VGND sg13g2_decap_4
XFILLER_3_161 VPWR VGND sg13g2_fill_1
X_3160_ _2752_ net896 net944 VPWR VGND sg13g2_nand2_1
Xhold1 mac1.sum_lvl1_ff\[41\] VPWR VGND net41 sg13g2_dlygate4sd3_1
X_3091_ _2683_ _2682_ _2673_ _2685_ VPWR VGND sg13g2_a21o_1
X_5801_ net811 net827 net780 _2507_ VPWR VGND sg13g2_mux2_1
X_3993_ _0836_ _0835_ _0126_ VPWR VGND sg13g2_xor2_1
X_5732_ net925 net907 net775 _2440_ VPWR VGND sg13g2_mux2_1
X_5663_ _2372_ _2367_ _2371_ VPWR VGND sg13g2_xnor2_1
X_5594_ mac2.total_sum\[4\] mac1.total_sum\[4\] _2316_ VPWR VGND sg13g2_xor2_1
X_4614_ _1429_ net827 net878 VPWR VGND sg13g2_nand2_1
Xhold401 DP_3.matrix\[8\] VPWR VGND net441 sg13g2_dlygate4sd3_1
X_4545_ _1358_ VPWR _1363_ VGND _1359_ _1361_ sg13g2_o21ai_1
Xhold445 _2159_ VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold412 _2255_ VPWR VGND net452 sg13g2_dlygate4sd3_1
Xhold423 _0042_ VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold434 mac2.sum_lvl3_ff\[20\] VPWR VGND net474 sg13g2_dlygate4sd3_1
X_4476_ _1281_ _1275_ _1283_ _1300_ VPWR VGND sg13g2_a21o_1
Xhold478 mac1.sum_lvl3_ff\[7\] VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold456 _0009_ VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold467 _2215_ VPWR VGND net507 sg13g2_dlygate4sd3_1
X_3427_ _0290_ _0269_ _0291_ VPWR VGND sg13g2_xor2_1
Xhold489 mac1.sum_lvl2_ff\[5\] VPWR VGND net529 sg13g2_dlygate4sd3_1
X_6215_ net1022 VGND VPWR net172 mac1.sum_lvl2_ff\[42\] clknet_leaf_66_clk sg13g2_dfrbpq_1
Xfanout903 net904 net903 VPWR VGND sg13g2_buf_2
Xfanout914 net915 net914 VPWR VGND sg13g2_buf_8
Xfanout925 net387 net925 VPWR VGND sg13g2_buf_8
X_6146_ net1075 VGND VPWR _0251_ DP_4.matrix\[7\] clknet_leaf_26_clk sg13g2_dfrbpq_2
Xfanout958 net959 net958 VPWR VGND sg13g2_buf_8
Xfanout936 net443 net936 VPWR VGND sg13g2_buf_1
Xfanout947 net948 net947 VPWR VGND sg13g2_buf_1
X_3358_ _2944_ _2939_ _2942_ VPWR VGND sg13g2_xnor2_1
Xfanout969 net970 net969 VPWR VGND sg13g2_buf_2
X_6077_ net1086 VGND VPWR _0204_ DP_2.matrix\[36\] clknet_leaf_50_clk sg13g2_dfrbpq_2
X_3289_ VGND VPWR _2843_ _2845_ _2878_ _2877_ sg13g2_a21oi_1
XFILLER_26_511 VPWR VGND sg13g2_fill_2
X_5028_ _1826_ net846 net787 VPWR VGND sg13g2_nand2_1
XFILLER_14_728 VPWR VGND sg13g2_fill_2
XFILLER_22_783 VPWR VGND sg13g2_fill_2
XFILLER_10_978 VPWR VGND sg13g2_decap_8
XFILLER_5_426 VPWR VGND sg13g2_fill_1
XFILLER_49_614 VPWR VGND sg13g2_decap_8
XFILLER_44_374 VPWR VGND sg13g2_fill_1
XFILLER_8_220 VPWR VGND sg13g2_fill_1
XFILLER_9_787 VPWR VGND sg13g2_fill_1
XFILLER_40_591 VPWR VGND sg13g2_fill_2
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_4330_ _1112_ VPWR _1159_ VGND _1052_ _1113_ sg13g2_o21ai_1
X_4261_ _1091_ net810 net864 VPWR VGND sg13g2_nand2_1
X_3212_ _2803_ _2797_ _2801_ VPWR VGND sg13g2_xnor2_1
X_6000_ net1070 VGND VPWR _0115_ mac1.products_ff\[9\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_4192_ _1024_ net868 net807 VPWR VGND sg13g2_nand2_1
X_3143_ _2735_ net954 net887 VPWR VGND sg13g2_nand2_1
X_3074_ _2668_ net956 net890 VPWR VGND sg13g2_nand2_1
XFILLER_39_179 VPWR VGND sg13g2_fill_1
XFILLER_39_1014 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_4
XFILLER_35_385 VPWR VGND sg13g2_fill_1
X_3976_ _0820_ net1008 net919 net960 net917 VPWR VGND sg13g2_a22oi_1
XFILLER_23_558 VPWR VGND sg13g2_decap_4
X_5715_ _2423_ _2421_ _2422_ _2420_ net770 VPWR VGND sg13g2_a22oi_1
X_5646_ _2354_ VPWR _2357_ VGND _2353_ _2355_ sg13g2_o21ai_1
Xhold220 mac1.sum_lvl2_ff\[41\] VPWR VGND net260 sg13g2_dlygate4sd3_1
X_5577_ _0054_ _2302_ net368 VPWR VGND sg13g2_xnor2_1
Xhold242 DP_4.matrix\[72\] VPWR VGND net282 sg13g2_dlygate4sd3_1
Xhold253 mac1.sum_lvl3_ff\[9\] VPWR VGND net293 sg13g2_dlygate4sd3_1
X_4528_ _1348_ net884 net829 _0084_ VPWR VGND sg13g2_and3_2
Xhold231 DP_3.matrix\[76\] VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold275 DP_4.matrix\[78\] VPWR VGND net315 sg13g2_dlygate4sd3_1
X_4459_ _1282_ _1274_ _1284_ VPWR VGND sg13g2_xor2_1
Xhold264 DP_1.matrix\[73\] VPWR VGND net304 sg13g2_dlygate4sd3_1
Xhold286 DP_1.matrix\[75\] VPWR VGND net326 sg13g2_dlygate4sd3_1
Xhold297 DP_4.matrix\[36\] VPWR VGND net337 sg13g2_dlygate4sd3_1
Xfanout766 _2454_ net766 VPWR VGND sg13g2_buf_8
Xfanout755 net756 net755 VPWR VGND sg13g2_buf_8
Xfanout788 net296 net788 VPWR VGND sg13g2_buf_8
Xfanout777 net778 net777 VPWR VGND sg13g2_buf_8
Xfanout799 net800 net799 VPWR VGND sg13g2_buf_2
X_6129_ net1054 VGND VPWR _0239_ DP_3.matrix\[75\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_39_680 VPWR VGND sg13g2_fill_1
XFILLER_27_875 VPWR VGND sg13g2_decap_8
XFILLER_42_889 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_fill_1
XFILLER_2_985 VPWR VGND sg13g2_decap_8
XFILLER_49_499 VPWR VGND sg13g2_fill_1
X_3830_ _0674_ _0675_ _0638_ _0678_ VPWR VGND sg13g2_nand3_1
X_3761_ net977 net924 _0074_ VPWR VGND sg13g2_and2_1
X_5500_ _2244_ mac2.sum_lvl2_ff\[33\] mac2.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_9_540 VPWR VGND sg13g2_fill_1
X_6480_ net1017 VGND VPWR net439 mac2.total_sum\[8\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3692_ _0549_ _0542_ _0548_ VPWR VGND sg13g2_xnor2_1
X_5431_ VGND VPWR _2184_ _2185_ _2191_ _2186_ sg13g2_a21oi_1
X_5362_ _2134_ VPWR _2137_ VGND _2133_ _2135_ sg13g2_o21ai_1
X_4313_ _1142_ net999 net817 net855 net814 VPWR VGND sg13g2_a22oi_1
X_5293_ _2083_ _2077_ _2082_ VPWR VGND sg13g2_xnor2_1
X_4244_ _1072_ _1071_ _1054_ _1075_ VPWR VGND sg13g2_a21o_1
X_4175_ _1008_ net867 net811 VPWR VGND sg13g2_nand2_1
X_3126_ _2707_ VPWR _2719_ VGND _2715_ _2717_ sg13g2_o21ai_1
X_3057_ _2641_ _2649_ _2651_ _2652_ VPWR VGND sg13g2_or3_1
XFILLER_24_812 VPWR VGND sg13g2_fill_2
XFILLER_36_683 VPWR VGND sg13g2_fill_1
XFILLER_36_694 VPWR VGND sg13g2_decap_8
X_3959_ _0803_ net971 net908 VPWR VGND sg13g2_nand2_1
XFILLER_13_1017 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_5629_ _2343_ _2336_ _2341_ VPWR VGND sg13g2_nand2_1
XFILLER_47_904 VPWR VGND sg13g2_decap_8
XFILLER_15_856 VPWR VGND sg13g2_fill_2
XFILLER_6_587 VPWR VGND sg13g2_fill_2
X_5980_ net792 _0262_ VPWR VGND sg13g2_buf_1
X_4931_ _1733_ _1732_ _1725_ VPWR VGND sg13g2_nand2b_1
X_4862_ _1670_ net877 net996 VPWR VGND sg13g2_nand2_1
XFILLER_33_664 VPWR VGND sg13g2_fill_1
X_3813_ _0659_ _0656_ _0661_ VPWR VGND sg13g2_xor2_1
X_4793_ _1484_ _1529_ _1483_ _1604_ VPWR VGND _1569_ sg13g2_nand4_1
X_3744_ _0597_ _0596_ _0599_ VPWR VGND sg13g2_xor2_1
X_3675_ _0498_ _0531_ _0496_ _0533_ VPWR VGND sg13g2_nand3_1
X_6463_ net1035 VGND VPWR _0045_ mac2.sum_lvl3_ff\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5414_ _2177_ _2172_ _2174_ VPWR VGND sg13g2_nand2_1
X_6394_ net1076 VGND VPWR net248 mac2.sum_lvl1_ff\[7\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5345_ _2123_ _2116_ _2121_ VPWR VGND sg13g2_nand2_1
X_5276_ _2042_ VPWR _2067_ VGND _2014_ _2040_ sg13g2_o21ai_1
X_4227_ _1057_ _1024_ _1058_ VPWR VGND sg13g2_xor2_1
XFILLER_29_937 VPWR VGND sg13g2_decap_8
XFILLER_44_907 VPWR VGND sg13g2_decap_8
X_4158_ net819 net813 net867 net865 _0992_ VPWR VGND sg13g2_and4_1
X_3109_ _2683_ _2673_ _2681_ _2702_ VPWR VGND sg13g2_a21o_1
X_4089_ VGND VPWR _0929_ _0930_ _0928_ _0870_ sg13g2_a21oi_2
XFILLER_24_620 VPWR VGND sg13g2_fill_2
XFILLER_12_815 VPWR VGND sg13g2_fill_2
XFILLER_8_808 VPWR VGND sg13g2_fill_1
XFILLER_3_524 VPWR VGND sg13g2_fill_1
XFILLER_3_513 VPWR VGND sg13g2_fill_1
XFILLER_11_85 VPWR VGND sg13g2_fill_2
XFILLER_3_579 VPWR VGND sg13g2_fill_2
XFILLER_19_403 VPWR VGND sg13g2_fill_2
XFILLER_35_929 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_43_962 VPWR VGND sg13g2_decap_8
XFILLER_15_664 VPWR VGND sg13g2_decap_8
Xinput13 uio_in[4] net13 VPWR VGND sg13g2_buf_1
X_3460_ _0322_ _0289_ _0323_ VPWR VGND sg13g2_xor2_1
X_3391_ net937 net932 net989 net987 _2972_ VPWR VGND sg13g2_and4_1
X_5130_ _1926_ _1921_ _1925_ VPWR VGND sg13g2_nand2_1
X_5061_ _1858_ net850 net781 VPWR VGND sg13g2_nand2_1
X_4012_ _0855_ net961 net914 net963 net913 VPWR VGND sg13g2_a22oi_1
XFILLER_38_745 VPWR VGND sg13g2_decap_4
X_5963_ net853 _0237_ VPWR VGND sg13g2_buf_1
X_4914_ _1716_ net289 _0090_ VPWR VGND sg13g2_nor2_1
XFILLER_34_940 VPWR VGND sg13g2_decap_8
X_5894_ _2574_ net829 net758 VPWR VGND sg13g2_nand2_1
X_4845_ VGND VPWR _1609_ _1614_ _1654_ _1626_ sg13g2_a21oi_1
X_4776_ _1587_ net823 net872 VPWR VGND sg13g2_nand2_1
XFILLER_20_177 VPWR VGND sg13g2_fill_2
X_3727_ _0583_ _0582_ _0565_ VPWR VGND sg13g2_nand2b_1
X_3658_ VPWR _0516_ _0515_ VGND sg13g2_inv_1
X_6446_ net1070 VGND VPWR net246 mac2.sum_lvl2_ff\[25\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_3589_ _0449_ _0398_ _0446_ VPWR VGND sg13g2_xnor2_1
X_6377_ net1035 VGND VPWR _0156_ mac2.products_ff\[142\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5328_ VGND VPWR _2105_ _2107_ _2110_ _2109_ sg13g2_a21oi_1
X_5259_ _2051_ _2036_ _2050_ VPWR VGND sg13g2_nand2_1
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_44_748 VPWR VGND sg13g2_fill_1
XFILLER_44_726 VPWR VGND sg13g2_fill_2
XFILLER_43_203 VPWR VGND sg13g2_fill_1
XFILLER_19_1001 VPWR VGND sg13g2_decap_8
XFILLER_25_973 VPWR VGND sg13g2_decap_8
XFILLER_12_645 VPWR VGND sg13g2_decap_8
XFILLER_11_155 VPWR VGND sg13g2_decap_8
XFILLER_40_976 VPWR VGND sg13g2_decap_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_520 VPWR VGND sg13g2_fill_2
XFILLER_19_299 VPWR VGND sg13g2_fill_1
XFILLER_16_984 VPWR VGND sg13g2_decap_8
XFILLER_31_976 VPWR VGND sg13g2_decap_8
X_4630_ _1445_ _1416_ _1444_ VPWR VGND sg13g2_nand2b_1
X_6300_ net1019 VGND VPWR _0015_ mac1.sum_lvl3_ff\[9\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4561_ _1378_ net878 net834 net880 net830 VPWR VGND sg13g2_a22oi_1
X_4492_ _1314_ _1300_ _1316_ VPWR VGND sg13g2_xor2_1
XFILLER_7_693 VPWR VGND sg13g2_decap_4
X_3512_ _0371_ _0372_ _0354_ _0374_ VPWR VGND sg13g2_nand3_1
X_3443_ _0305_ _0304_ _0287_ _0307_ VPWR VGND sg13g2_a21o_1
X_6231_ net1049 VGND VPWR net95 mac2.sum_lvl2_ff\[42\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_6162_ net1061 VGND VPWR _0267_ DP_4.matrix\[79\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3374_ _2959_ _2946_ _2958_ VPWR VGND sg13g2_xnor2_1
X_5113_ _1908_ _1904_ _1909_ VPWR VGND sg13g2_xor2_1
X_6093_ net1042 VGND VPWR _0215_ DP_2.matrix\[75\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5044_ _1830_ VPWR _1842_ VGND _1838_ _1840_ sg13g2_o21ai_1
XFILLER_38_597 VPWR VGND sg13g2_decap_8
X_5946_ net277 _0212_ VPWR VGND sg13g2_buf_1
X_5877_ _2471_ _2460_ _2563_ VPWR VGND sg13g2_xor2_1
X_4828_ _1637_ DP_4.matrix\[5\] net1001 VPWR VGND sg13g2_nand2_2
XFILLER_22_976 VPWR VGND sg13g2_decap_8
XFILLER_21_497 VPWR VGND sg13g2_fill_2
X_4759_ _1570_ _1569_ _0148_ VPWR VGND sg13g2_xor2_1
X_6429_ net1076 VGND VPWR net140 mac2.sum_lvl2_ff\[5\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_44_512 VPWR VGND sg13g2_fill_1
XFILLER_1_1018 VPWR VGND sg13g2_decap_8
XFILLER_32_718 VPWR VGND sg13g2_decap_4
XFILLER_13_954 VPWR VGND sg13g2_decap_8
XFILLER_12_486 VPWR VGND sg13g2_fill_2
XFILLER_8_468 VPWR VGND sg13g2_fill_2
XFILLER_3_195 VPWR VGND sg13g2_fill_1
X_3090_ _2682_ _2683_ _2673_ _2684_ VPWR VGND sg13g2_nand3_1
Xhold2 mac2.sum_lvl1_ff\[81\] VPWR VGND net42 sg13g2_dlygate4sd3_1
XFILLER_48_884 VPWR VGND sg13g2_decap_8
X_3992_ _0836_ _0793_ _0796_ VPWR VGND sg13g2_nand2_1
X_5800_ _2501_ _2505_ _2506_ VPWR VGND sg13g2_nor2b_1
X_5731_ _2439_ _2436_ _2438_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_291 VPWR VGND sg13g2_fill_1
X_5662_ _2371_ DP_1.I_range.out_data\[2\] VPWR VGND DP_1.Q_range.out_data\[2\] sg13g2_nand2b_2
X_5593_ mac1.total_sum\[4\] mac2.total_sum\[4\] _2315_ VPWR VGND sg13g2_and2_1
X_4613_ _1399_ VPWR _1428_ VGND _1397_ _1400_ sg13g2_o21ai_1
XFILLER_8_980 VPWR VGND sg13g2_decap_8
Xhold402 DP_2.matrix\[37\] VPWR VGND net442 sg13g2_dlygate4sd3_1
X_4544_ _1358_ _1359_ _1361_ _1362_ VPWR VGND sg13g2_nor3_1
Xhold413 _0056_ VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold435 _0055_ VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold424 DP_2.matrix\[43\] VPWR VGND net464 sg13g2_dlygate4sd3_1
Xhold457 DP_3.matrix\[41\] VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold446 _0028_ VPWR VGND net486 sg13g2_dlygate4sd3_1
X_6214_ net1024 VGND VPWR net87 mac1.sum_lvl2_ff\[41\] clknet_leaf_65_clk sg13g2_dfrbpq_1
Xhold468 _0046_ VPWR VGND net508 sg13g2_dlygate4sd3_1
X_4475_ _1289_ _1269_ _1288_ _1299_ VPWR VGND sg13g2_a21o_1
X_3426_ _0290_ net990 net929 VPWR VGND sg13g2_nand2_1
Xfanout915 net504 net915 VPWR VGND sg13g2_buf_2
Xfanout904 net905 net904 VPWR VGND sg13g2_buf_2
Xhold479 _2161_ VPWR VGND net519 sg13g2_dlygate4sd3_1
X_6145_ net1075 VGND VPWR _0250_ DP_4.matrix\[6\] clknet_leaf_26_clk sg13g2_dfrbpq_2
Xfanout948 net336 net948 VPWR VGND sg13g2_buf_1
Xfanout937 net940 net937 VPWR VGND sg13g2_buf_8
X_3357_ _2943_ _2942_ _2939_ VPWR VGND sg13g2_nand2b_1
Xfanout926 net414 net926 VPWR VGND sg13g2_buf_8
Xfanout959 net299 net959 VPWR VGND sg13g2_buf_8
X_6076_ net1017 VGND VPWR _0104_ mac1.products_ff\[145\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3288_ _2875_ _2853_ _2877_ VPWR VGND sg13g2_xor2_1
X_5027_ _1825_ net850 net785 VPWR VGND sg13g2_nand2_1
XFILLER_39_895 VPWR VGND sg13g2_decap_8
X_5929_ net961 _0187_ VPWR VGND sg13g2_buf_1
XFILLER_16_1026 VPWR VGND sg13g2_fill_2
XFILLER_21_272 VPWR VGND sg13g2_fill_2
XFILLER_10_957 VPWR VGND sg13g2_decap_8
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_44_93 VPWR VGND sg13g2_fill_2
XFILLER_32_559 VPWR VGND sg13g2_decap_4
XFILLER_12_272 VPWR VGND sg13g2_fill_1
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_4260_ _1090_ net868 net805 VPWR VGND sg13g2_nand2_1
X_3211_ _2802_ _2797_ _2801_ VPWR VGND sg13g2_nand2_1
X_4191_ _1023_ net871 net806 VPWR VGND sg13g2_nand2_1
X_3142_ _2734_ net959 net1003 VPWR VGND sg13g2_nand2_1
X_3073_ _2650_ VPWR _2667_ VGND _2641_ _2651_ sg13g2_o21ai_1
X_3975_ net919 net917 net960 net1008 _0819_ VPWR VGND sg13g2_and4_1
X_5714_ net770 VPWR _2422_ VGND net918 net774 sg13g2_o21ai_1
X_5645_ net23 _2353_ _2356_ VPWR VGND sg13g2_xnor2_1
Xhold210 mac2.sum_lvl1_ff\[87\] VPWR VGND net250 sg13g2_dlygate4sd3_1
X_5576_ _2303_ mac2.sum_lvl3_ff\[35\] net367 VPWR VGND sg13g2_xnor2_1
Xhold232 DP_4.matrix\[80\] VPWR VGND net272 sg13g2_dlygate4sd3_1
Xhold221 mac2.products_ff\[13\] VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold243 mac1.sum_lvl3_ff\[0\] VPWR VGND net283 sg13g2_dlygate4sd3_1
X_4527_ net886 net833 _0084_ VPWR VGND sg13g2_and2_1
XFILLER_46_1008 VPWR VGND sg13g2_decap_8
Xhold276 DP_3.matrix\[80\] VPWR VGND net316 sg13g2_dlygate4sd3_1
X_4458_ _1282_ _1274_ _1283_ VPWR VGND sg13g2_nor2b_1
Xhold254 _2170_ VPWR VGND net294 sg13g2_dlygate4sd3_1
Xhold265 mac2.sum_lvl3_ff\[0\] VPWR VGND net305 sg13g2_dlygate4sd3_1
Xhold287 DP_3.matrix\[38\] VPWR VGND net327 sg13g2_dlygate4sd3_1
X_3409_ net937 net936 net987 net985 _0274_ VPWR VGND sg13g2_and4_1
Xhold298 mac2.sum_lvl3_ff\[9\] VPWR VGND net338 sg13g2_dlygate4sd3_1
Xfanout756 net757 net756 VPWR VGND sg13g2_buf_8
X_6128_ net1056 VGND VPWR _0238_ DP_3.matrix\[74\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4389_ _1214_ _1206_ _1216_ VPWR VGND sg13g2_xor2_1
Xfanout767 net769 net767 VPWR VGND sg13g2_buf_8
Xfanout789 net790 net789 VPWR VGND sg13g2_buf_8
Xfanout778 _2449_ net778 VPWR VGND sg13g2_buf_1
X_6059_ net1041 VGND VPWR _0192_ DP_1.matrix\[76\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_14_548 VPWR VGND sg13g2_fill_2
XFILLER_42_868 VPWR VGND sg13g2_decap_8
XFILLER_22_592 VPWR VGND sg13g2_fill_2
XFILLER_2_964 VPWR VGND sg13g2_decap_8
XFILLER_7_1013 VPWR VGND sg13g2_decap_8
XFILLER_1_463 VPWR VGND sg13g2_fill_2
XFILLER_49_456 VPWR VGND sg13g2_fill_1
XFILLER_37_607 VPWR VGND sg13g2_decap_8
XFILLER_37_618 VPWR VGND sg13g2_fill_1
XFILLER_44_161 VPWR VGND sg13g2_fill_1
XFILLER_18_898 VPWR VGND sg13g2_decap_8
XFILLER_32_345 VPWR VGND sg13g2_fill_1
X_3760_ _0111_ _0606_ _0613_ VPWR VGND sg13g2_xnor2_1
X_5430_ net373 mac1.sum_lvl3_ff\[34\] _2190_ VPWR VGND sg13g2_xor2_1
X_3691_ _0548_ _0543_ _0546_ VPWR VGND sg13g2_xnor2_1
X_5361_ _0005_ _2133_ net469 VPWR VGND sg13g2_xnor2_1
X_5292_ _2082_ _2068_ _2081_ VPWR VGND sg13g2_xnor2_1
X_4312_ net814 net855 net817 _1141_ VPWR VGND net999 sg13g2_nand4_1
X_4243_ VGND VPWR _1071_ _1072_ _1074_ _1054_ sg13g2_a21oi_1
X_4174_ _0993_ VPWR _1007_ VGND _0991_ _0994_ sg13g2_o21ai_1
X_3125_ _2707_ _2715_ _2717_ _2718_ VPWR VGND sg13g2_or3_1
X_3056_ VGND VPWR _2647_ _2648_ _2651_ _2642_ sg13g2_a21oi_1
XFILLER_27_139 VPWR VGND sg13g2_fill_2
XFILLER_24_868 VPWR VGND sg13g2_fill_1
X_3958_ _0802_ net971 net906 VPWR VGND sg13g2_nand2_1
X_3889_ _0735_ _0728_ _0733_ _0734_ VPWR VGND sg13g2_and3_1
X_5628_ net20 _2341_ _2342_ VPWR VGND sg13g2_xnor2_1
X_5559_ _2278_ _2282_ _2288_ _2289_ VPWR VGND sg13g2_nor3_1
XFILLER_15_879 VPWR VGND sg13g2_fill_2
XFILLER_14_367 VPWR VGND sg13g2_fill_2
XFILLER_10_584 VPWR VGND sg13g2_decap_4
XFILLER_41_94 VPWR VGND sg13g2_decap_4
XFILLER_29_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_271 VPWR VGND sg13g2_fill_2
XFILLER_38_949 VPWR VGND sg13g2_decap_8
X_4930_ _1730_ _1731_ _1732_ VPWR VGND sg13g2_nor2b_1
X_4861_ _1645_ VPWR _1669_ VGND _1642_ _1646_ sg13g2_o21ai_1
XFILLER_17_183 VPWR VGND sg13g2_fill_2
XFILLER_36_1018 VPWR VGND sg13g2_decap_8
X_3812_ _0660_ _0659_ _0656_ VPWR VGND sg13g2_nand2b_1
XFILLER_33_698 VPWR VGND sg13g2_decap_4
X_4792_ _1601_ _1602_ _1603_ VPWR VGND sg13g2_nor2b_1
X_3743_ _0598_ _0596_ _0597_ VPWR VGND sg13g2_nand2_1
X_3674_ VGND VPWR _0496_ _0498_ _0532_ _0531_ sg13g2_a21oi_1
X_6462_ net1049 VGND VPWR net527 mac2.sum_lvl3_ff\[6\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5413_ _2176_ mac1.sum_lvl3_ff\[31\] net393 VPWR VGND sg13g2_xnor2_1
X_6393_ net1076 VGND VPWR net254 mac2.sum_lvl1_ff\[6\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5344_ _0002_ _2121_ _2122_ VPWR VGND sg13g2_xnor2_1
X_5275_ _2066_ _2061_ _2064_ VPWR VGND sg13g2_xnor2_1
X_4226_ _1057_ net866 net810 VPWR VGND sg13g2_nand2_1
XFILLER_29_916 VPWR VGND sg13g2_decap_8
X_4157_ _0991_ net869 net811 VPWR VGND sg13g2_nand2_1
X_3108_ _2701_ _2695_ _2699_ VPWR VGND sg13g2_xnor2_1
X_4088_ _0898_ VPWR _0929_ VGND _0868_ _0897_ sg13g2_o21ai_1
X_3039_ _2633_ _2615_ _0068_ VPWR VGND sg13g2_xor2_1
XFILLER_37_993 VPWR VGND sg13g2_decap_8
XFILLER_23_153 VPWR VGND sg13g2_fill_1
XFILLER_47_746 VPWR VGND sg13g2_fill_2
XFILLER_35_908 VPWR VGND sg13g2_decap_8
XFILLER_28_993 VPWR VGND sg13g2_decap_8
XFILLER_43_941 VPWR VGND sg13g2_decap_8
Xinput14 uio_in[5] net14 VPWR VGND sg13g2_buf_1
XFILLER_10_370 VPWR VGND sg13g2_fill_2
X_3390_ _2971_ net991 net930 VPWR VGND sg13g2_nand2_1
X_5060_ _1857_ net854 net994 VPWR VGND sg13g2_nand2_1
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
X_4011_ net914 net912 net963 net961 _0854_ VPWR VGND sg13g2_and4_1
XFILLER_37_212 VPWR VGND sg13g2_fill_1
XFILLER_38_724 VPWR VGND sg13g2_decap_4
XFILLER_26_908 VPWR VGND sg13g2_fill_2
XFILLER_26_919 VPWR VGND sg13g2_decap_4
X_5962_ net279 _0236_ VPWR VGND sg13g2_buf_1
X_4913_ _1717_ net796 net279 net853 net800 VPWR VGND sg13g2_a22oi_1
XFILLER_33_451 VPWR VGND sg13g2_fill_1
XFILLER_34_996 VPWR VGND sg13g2_decap_8
X_5893_ _2505_ _2501_ _2573_ VPWR VGND sg13g2_xor2_1
X_4844_ _1651_ _1639_ _1653_ VPWR VGND sg13g2_xor2_1
XFILLER_21_635 VPWR VGND sg13g2_decap_4
X_4775_ _1586_ net877 net822 VPWR VGND sg13g2_nand2_1
XFILLER_21_657 VPWR VGND sg13g2_decap_8
X_3726_ _0582_ _0566_ _0580_ VPWR VGND sg13g2_xnor2_1
X_3657_ _0478_ VPWR _0515_ VGND _0475_ _0479_ sg13g2_o21ai_1
X_6445_ net1076 VGND VPWR net72 mac2.sum_lvl2_ff\[24\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3588_ _0398_ _0446_ _0448_ VPWR VGND sg13g2_and2_1
X_6376_ net1036 VGND VPWR _0149_ mac2.products_ff\[141\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5327_ _2109_ mac1.sum_lvl2_ff\[27\] mac1.sum_lvl2_ff\[8\] VPWR VGND sg13g2_xnor2_1
X_5258_ _2050_ _2022_ _2048_ VPWR VGND sg13g2_xnor2_1
X_5189_ _1982_ _1979_ _1983_ VPWR VGND sg13g2_xor2_1
X_4209_ _1039_ _1040_ _1022_ _1041_ VPWR VGND sg13g2_nand3_1
XFILLER_44_705 VPWR VGND sg13g2_fill_1
XFILLER_25_941 VPWR VGND sg13g2_fill_2
XFILLER_25_952 VPWR VGND sg13g2_decap_8
XFILLER_11_123 VPWR VGND sg13g2_fill_1
XFILLER_40_955 VPWR VGND sg13g2_decap_8
XFILLER_12_668 VPWR VGND sg13g2_fill_1
XFILLER_8_639 VPWR VGND sg13g2_fill_1
XFILLER_7_127 VPWR VGND sg13g2_fill_1
XFILLER_4_878 VPWR VGND sg13g2_fill_1
XFILLER_4_889 VPWR VGND sg13g2_decap_8
XFILLER_26_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_278 VPWR VGND sg13g2_decap_8
XFILLER_16_963 VPWR VGND sg13g2_decap_8
XFILLER_31_955 VPWR VGND sg13g2_decap_8
X_4560_ net830 net880 net834 _1377_ VPWR VGND net878 sg13g2_nand4_1
X_4491_ _1315_ _1300_ _1314_ VPWR VGND sg13g2_nand2_1
X_3511_ _0373_ _0354_ _0371_ _0372_ VPWR VGND sg13g2_and3_1
X_3442_ _0304_ _0305_ _0287_ _0306_ VPWR VGND sg13g2_nand3_1
X_6230_ net1051 VGND VPWR net84 mac2.sum_lvl2_ff\[41\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6161_ net1055 VGND VPWR _0266_ DP_4.matrix\[78\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3373_ _2958_ _2955_ _2957_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_2 VPWR VGND sg13g2_fill_1
X_5112_ _1908_ _1858_ _1906_ VPWR VGND sg13g2_xnor2_1
X_6092_ net1063 VGND VPWR _0214_ DP_2.matrix\[74\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_26_0 VPWR VGND sg13g2_fill_2
XFILLER_38_521 VPWR VGND sg13g2_fill_1
X_5043_ _1830_ _1838_ _1840_ _1841_ VPWR VGND sg13g2_or3_1
X_5945_ net906 _0211_ VPWR VGND sg13g2_buf_1
X_5876_ _2562_ VPWR _0222_ VGND net758 _2561_ sg13g2_o21ai_1
X_4827_ _1636_ net1002 net824 net872 DP_4.matrix\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_22_955 VPWR VGND sg13g2_decap_8
XFILLER_21_465 VPWR VGND sg13g2_fill_1
X_4758_ _1570_ _1527_ _1530_ VPWR VGND sg13g2_nand2_1
X_3709_ _0556_ _0536_ _0555_ _0565_ VPWR VGND sg13g2_a21o_1
X_4689_ _1498_ _1500_ _1501_ _1502_ VPWR VGND sg13g2_nor3_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_1017 VPWR VGND sg13g2_decap_8
X_6428_ net1073 VGND VPWR net90 mac2.sum_lvl2_ff\[4\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_6359_ net1072 VGND VPWR _0083_ mac2.products_ff\[72\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_17_30 VPWR VGND sg13g2_fill_1
XFILLER_29_565 VPWR VGND sg13g2_fill_2
XFILLER_13_922 VPWR VGND sg13g2_fill_2
XFILLER_9_915 VPWR VGND sg13g2_fill_2
XFILLER_9_959 VPWR VGND sg13g2_decap_8
Xhold3 mac1.products_ff\[144\] VPWR VGND net43 sg13g2_dlygate4sd3_1
XFILLER_0_892 VPWR VGND sg13g2_decap_8
XFILLER_48_863 VPWR VGND sg13g2_decap_8
X_3991_ _0832_ _0834_ _0835_ VPWR VGND sg13g2_nor2_1
X_5730_ _2438_ net772 _2437_ net764 net280 VPWR VGND sg13g2_a22oi_1
X_5661_ _2367_ net776 _2370_ VPWR VGND sg13g2_nor2_2
X_5592_ _2312_ VPWR _2314_ VGND _2311_ _2313_ sg13g2_o21ai_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
X_4612_ _1427_ _1422_ _1425_ VPWR VGND sg13g2_xnor2_1
X_4543_ _1361_ net880 net834 net882 net829 VPWR VGND sg13g2_a22oi_1
Xhold425 DP_4.matrix\[43\] VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold436 DP_4.matrix\[8\] VPWR VGND net476 sg13g2_dlygate4sd3_1
XFILLER_7_480 VPWR VGND sg13g2_fill_1
Xhold403 DP_2.matrix\[1\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold414 mac2.sum_lvl3_ff\[4\] VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold469 DP_1.matrix\[3\] VPWR VGND net509 sg13g2_dlygate4sd3_1
X_6213_ net1039 VGND VPWR net115 mac1.sum_lvl2_ff\[40\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xhold447 mac2.sum_lvl3_ff\[3\] VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold458 DP_3.matrix\[2\] VPWR VGND net498 sg13g2_dlygate4sd3_1
X_4474_ _1297_ _1293_ _0130_ VPWR VGND sg13g2_xor2_1
Xfanout905 DP_2.matrix\[72\] net905 VPWR VGND sg13g2_buf_2
Xfanout916 net335 net916 VPWR VGND sg13g2_buf_8
X_3425_ _0289_ net990 net928 VPWR VGND sg13g2_nand2_1
X_6144_ net1075 VGND VPWR _0249_ DP_4.matrix\[5\] clknet_leaf_26_clk sg13g2_dfrbpq_2
Xfanout949 net951 net949 VPWR VGND sg13g2_buf_8
Xfanout938 net939 net938 VPWR VGND sg13g2_buf_2
X_3356_ _2941_ _2916_ _2942_ VPWR VGND sg13g2_xor2_1
Xfanout927 net422 net927 VPWR VGND sg13g2_buf_8
X_3287_ _2875_ _2853_ _2876_ VPWR VGND sg13g2_nor2b_1
X_6075_ net1065 VGND VPWR _0203_ DP_2.matrix\[7\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_5026_ _1805_ _1795_ _1803_ _1824_ VPWR VGND sg13g2_a21o_1
XFILLER_26_513 VPWR VGND sg13g2_fill_1
XFILLER_39_874 VPWR VGND sg13g2_decap_8
XFILLER_41_505 VPWR VGND sg13g2_decap_4
X_5928_ net963 _0186_ VPWR VGND sg13g2_buf_1
XFILLER_16_1005 VPWR VGND sg13g2_decap_8
XFILLER_10_936 VPWR VGND sg13g2_decap_8
X_5859_ _2434_ _2430_ _2552_ VPWR VGND sg13g2_xor2_1
XFILLER_22_785 VPWR VGND sg13g2_fill_1
XFILLER_0_111 VPWR VGND sg13g2_fill_2
XFILLER_0_122 VPWR VGND sg13g2_fill_1
XFILLER_49_649 VPWR VGND sg13g2_decap_8
XFILLER_45_888 VPWR VGND sg13g2_decap_8
XFILLER_17_557 VPWR VGND sg13g2_decap_8
XFILLER_9_701 VPWR VGND sg13g2_fill_1
XFILLER_13_741 VPWR VGND sg13g2_fill_1
XFILLER_40_560 VPWR VGND sg13g2_fill_2
XFILLER_5_951 VPWR VGND sg13g2_decap_8
X_3210_ _2799_ _2800_ _2801_ VPWR VGND sg13g2_nor2_1
X_4190_ _1014_ VPWR _1022_ VGND _1006_ _1016_ sg13g2_o21ai_1
X_3141_ _2705_ VPWR _2733_ VGND _2703_ _2706_ sg13g2_o21ai_1
X_3072_ _2664_ _2663_ _2666_ VPWR VGND sg13g2_xor2_1
XFILLER_48_682 VPWR VGND sg13g2_fill_2
XFILLER_23_516 VPWR VGND sg13g2_fill_1
XFILLER_35_398 VPWR VGND sg13g2_fill_2
XFILLER_36_899 VPWR VGND sg13g2_decap_8
X_3974_ _0818_ net916 net1008 VPWR VGND sg13g2_nand2_1
X_5713_ _2421_ net902 net774 VPWR VGND sg13g2_nand2_1
X_5644_ mac2.total_sum\[14\] mac1.total_sum\[14\] _2356_ VPWR VGND sg13g2_xor2_1
Xhold200 mac1.products_ff\[76\] VPWR VGND net240 sg13g2_dlygate4sd3_1
Xhold211 mac2.sum_lvl2_ff\[43\] VPWR VGND net251 sg13g2_dlygate4sd3_1
X_5575_ _2299_ VPWR _2302_ VGND _2298_ _2300_ sg13g2_o21ai_1
Xhold233 DP_4.matrix\[44\] VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold222 mac2.products_ff\[14\] VPWR VGND net262 sg13g2_dlygate4sd3_1
X_4526_ _0133_ _1340_ _1347_ VPWR VGND sg13g2_xnor2_1
Xhold244 _0016_ VPWR VGND net284 sg13g2_dlygate4sd3_1
XFILLER_2_409 VPWR VGND sg13g2_fill_2
X_4457_ _1282_ _1275_ _1281_ VPWR VGND sg13g2_xnor2_1
Xhold277 mac1.sum_lvl3_ff\[5\] VPWR VGND net317 sg13g2_dlygate4sd3_1
Xhold266 _0048_ VPWR VGND net306 sg13g2_dlygate4sd3_1
Xhold255 _0031_ VPWR VGND net295 sg13g2_dlygate4sd3_1
Xhold288 DP_4.matrix\[39\] VPWR VGND net328 sg13g2_dlygate4sd3_1
X_3408_ _0273_ net989 net930 VPWR VGND sg13g2_nand2_1
Xhold299 _2279_ VPWR VGND net339 sg13g2_dlygate4sd3_1
X_6127_ net1080 VGND VPWR net98 mac1.sum_lvl1_ff\[10\] clknet_leaf_43_clk sg13g2_dfrbpq_1
Xfanout757 _2366_ net757 VPWR VGND sg13g2_buf_8
X_4388_ _1214_ _1206_ _1215_ VPWR VGND sg13g2_nor2b_1
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_8
X_3339_ _2926_ _2925_ _2898_ VPWR VGND sg13g2_nand2b_1
Xfanout779 _2448_ net779 VPWR VGND sg13g2_buf_8
XFILLER_45_107 VPWR VGND sg13g2_fill_1
X_6058_ net1022 VGND VPWR _0067_ mac1.products_ff\[139\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_39_671 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_65_clk clknet_4_0_0_clk clknet_leaf_65_clk VPWR VGND sg13g2_buf_8
X_5009_ _1806_ _1807_ _1789_ _1808_ VPWR VGND sg13g2_nand3_1
XFILLER_41_302 VPWR VGND sg13g2_fill_1
XFILLER_2_943 VPWR VGND sg13g2_decap_8
XFILLER_49_435 VPWR VGND sg13g2_fill_2
XFILLER_18_800 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_56_clk clknet_4_8_0_clk clknet_leaf_56_clk VPWR VGND sg13g2_buf_8
XFILLER_18_877 VPWR VGND sg13g2_fill_2
XFILLER_32_368 VPWR VGND sg13g2_fill_1
X_3690_ _0547_ _0546_ _0543_ VPWR VGND sg13g2_nand2b_1
X_5360_ net468 mac1.sum_lvl2_ff\[33\] _2136_ VPWR VGND sg13g2_xor2_1
X_5291_ _2081_ _2078_ _2080_ VPWR VGND sg13g2_xnor2_1
X_4311_ net817 net814 net855 net999 _1140_ VPWR VGND sg13g2_and4_1
X_4242_ _1071_ _1072_ _1054_ _1073_ VPWR VGND sg13g2_nand3_1
X_4173_ VGND VPWR _1006_ _1005_ _1003_ sg13g2_or2_1
X_3124_ VGND VPWR _2713_ _2714_ _2717_ _2708_ sg13g2_a21oi_1
X_3055_ _2647_ _2648_ _2642_ _2650_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_47_clk clknet_4_14_0_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
X_3957_ _0801_ net976 net1004 VPWR VGND sg13g2_nand2_1
X_3888_ _0729_ VPWR _0734_ VGND _0730_ _0732_ sg13g2_o21ai_1
X_5627_ VGND VPWR _2336_ _2338_ _2342_ _2335_ sg13g2_a21oi_1
X_5558_ _2288_ _2281_ _2286_ VPWR VGND sg13g2_nand2_1
X_4509_ _1306_ VPWR _1332_ VGND _1277_ _1304_ sg13g2_o21ai_1
X_5489_ _2230_ _2225_ _2229_ _2235_ VPWR VGND sg13g2_a21o_1
XFILLER_47_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_38_clk clknet_4_15_0_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_14_313 VPWR VGND sg13g2_fill_1
XFILLER_41_62 VPWR VGND sg13g2_decap_4
XFILLER_6_589 VPWR VGND sg13g2_fill_1
XFILLER_37_8 VPWR VGND sg13g2_fill_1
XFILLER_38_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_4_12_0_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_46_994 VPWR VGND sg13g2_decap_8
X_4860_ _1648_ _1641_ _1650_ _1668_ VPWR VGND sg13g2_a21o_1
X_3811_ _0658_ _0637_ _0659_ VPWR VGND sg13g2_xor2_1
X_4791_ _1564_ _1600_ _1562_ _1602_ VPWR VGND sg13g2_nand3_1
X_3742_ _0572_ VPWR _0597_ VGND _0544_ _0570_ sg13g2_o21ai_1
X_3673_ _0529_ _0506_ _0531_ VPWR VGND sg13g2_xor2_1
X_6461_ net1049 VGND VPWR net450 mac2.sum_lvl3_ff\[5\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5412_ mac1.sum_lvl3_ff\[31\] mac1.sum_lvl3_ff\[11\] _2175_ VPWR VGND sg13g2_nor2_1
X_6392_ net1073 VGND VPWR net122 mac2.sum_lvl1_ff\[5\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5343_ VGND VPWR _2116_ _2118_ _2122_ _2115_ sg13g2_a21oi_1
X_5274_ _2065_ _2064_ _2061_ VPWR VGND sg13g2_nand2b_1
X_4225_ _1056_ net866 net807 VPWR VGND sg13g2_nand2_1
X_4156_ VGND VPWR _0983_ _0986_ _0990_ _0984_ sg13g2_a21oi_1
X_3107_ _2695_ _2699_ _2700_ VPWR VGND sg13g2_and2_1
X_4087_ _0871_ _0927_ _0928_ VPWR VGND sg13g2_nor2b_1
X_3038_ _2615_ _2633_ _2634_ VPWR VGND sg13g2_and2_1
XFILLER_37_972 VPWR VGND sg13g2_decap_8
XFILLER_12_817 VPWR VGND sg13g2_fill_1
X_4989_ _1786_ _1785_ _1788_ VPWR VGND sg13g2_xor2_1
XFILLER_19_405 VPWR VGND sg13g2_fill_1
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_4_1017 VPWR VGND sg13g2_decap_8
XFILLER_43_920 VPWR VGND sg13g2_decap_8
XFILLER_28_972 VPWR VGND sg13g2_decap_8
XFILLER_43_997 VPWR VGND sg13g2_decap_8
XFILLER_30_636 VPWR VGND sg13g2_fill_2
Xheichips25_SDR_40 VPWR VGND uio_oe[7] sg13g2_tiehi
Xinput15 uio_in[6] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_887 VPWR VGND sg13g2_fill_2
XFILLER_42_1001 VPWR VGND sg13g2_decap_8
X_4010_ _0853_ net912 net961 VPWR VGND sg13g2_nand2_1
XFILLER_28_4 VPWR VGND sg13g2_fill_1
XFILLER_38_769 VPWR VGND sg13g2_decap_8
X_5961_ net856 _0235_ VPWR VGND sg13g2_buf_1
XFILLER_19_994 VPWR VGND sg13g2_decap_8
X_4912_ _1716_ net853 net796 _0089_ VPWR VGND sg13g2_and3_2
X_5892_ _0244_ net833 net758 VPWR VGND sg13g2_xnor2_1
XFILLER_34_975 VPWR VGND sg13g2_decap_8
X_4843_ VGND VPWR _1652_ _1651_ _1639_ sg13g2_or2_1
X_4774_ VGND VPWR net831 net872 _1585_ _1552_ sg13g2_a21oi_1
X_3725_ _0581_ _0566_ _0580_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_9_clk clknet_4_3_0_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_6444_ net1073 VGND VPWR net69 mac2.sum_lvl2_ff\[23\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3656_ _0514_ _0508_ _0513_ VPWR VGND sg13g2_xnor2_1
X_3587_ VGND VPWR _0447_ _0445_ _0399_ sg13g2_or2_1
X_6375_ net1036 VGND VPWR _0093_ mac2.products_ff\[140\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5326_ _2107_ _2108_ _0013_ VPWR VGND sg13g2_and2_1
X_5257_ _2049_ _2048_ _2022_ VPWR VGND sg13g2_nand2b_1
X_4208_ _1028_ VPWR _1040_ VGND _1036_ _1038_ sg13g2_o21ai_1
X_5188_ _1982_ _1957_ _1980_ VPWR VGND sg13g2_xnor2_1
X_4139_ _0977_ _0960_ _0976_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_728 VPWR VGND sg13g2_fill_1
XFILLER_43_238 VPWR VGND sg13g2_fill_2
XFILLER_40_934 VPWR VGND sg13g2_decap_8
XFILLER_11_168 VPWR VGND sg13g2_fill_1
XFILLER_47_522 VPWR VGND sg13g2_fill_1
XFILLER_35_706 VPWR VGND sg13g2_decap_4
XFILLER_47_588 VPWR VGND sg13g2_fill_2
XFILLER_47_566 VPWR VGND sg13g2_fill_2
XFILLER_47_94 VPWR VGND sg13g2_fill_2
XFILLER_34_205 VPWR VGND sg13g2_fill_1
XFILLER_16_920 VPWR VGND sg13g2_fill_2
XFILLER_15_430 VPWR VGND sg13g2_fill_2
XFILLER_43_794 VPWR VGND sg13g2_decap_4
XFILLER_31_934 VPWR VGND sg13g2_decap_8
XFILLER_42_260 VPWR VGND sg13g2_fill_1
X_3510_ _0360_ VPWR _0372_ VGND _0368_ _0370_ sg13g2_o21ai_1
X_4490_ _1314_ _1285_ _1312_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_150 VPWR VGND sg13g2_fill_2
X_3441_ _0293_ VPWR _0305_ VGND _0301_ _0303_ sg13g2_o21ai_1
X_6160_ net1060 VGND VPWR _0265_ DP_4.matrix\[77\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3372_ _2957_ _2940_ _2956_ VPWR VGND sg13g2_xnor2_1
X_5111_ VGND VPWR _1907_ _1905_ _1859_ sg13g2_or2_1
X_6091_ net1042 VGND VPWR _0099_ mac1.products_ff\[150\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5042_ VGND VPWR _1836_ _1837_ _1840_ _1831_ sg13g2_a21oi_1
X_5944_ net908 _0210_ VPWR VGND sg13g2_buf_1
X_5875_ _2562_ net882 net758 VPWR VGND sg13g2_nand2_1
X_4826_ VGND VPWR _1617_ _1622_ _1635_ _1624_ sg13g2_a21oi_1
XFILLER_21_499 VPWR VGND sg13g2_fill_1
X_4757_ _1566_ _1568_ _1569_ VPWR VGND sg13g2_nor2_1
X_3708_ _0564_ _0560_ _0108_ VPWR VGND sg13g2_xor2_1
X_4688_ _1501_ net877 net826 net823 net879 VPWR VGND sg13g2_a22oi_1
X_3639_ _0498_ _0471_ _0497_ VPWR VGND sg13g2_nand2_1
X_6427_ net1072 VGND VPWR net109 mac2.sum_lvl2_ff\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_1_805 VPWR VGND sg13g2_fill_2
X_6358_ net1072 VGND VPWR _0082_ mac2.products_ff\[71\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5309_ mac1.sum_lvl2_ff\[23\] mac1.sum_lvl2_ff\[4\] _2095_ VPWR VGND sg13g2_and2_1
X_6289_ net1046 VGND VPWR net226 mac1.sum_lvl3_ff\[34\] clknet_leaf_10_clk sg13g2_dfrbpq_2
XFILLER_13_901 VPWR VGND sg13g2_decap_4
XFILLER_40_731 VPWR VGND sg13g2_decap_4
XFILLER_40_742 VPWR VGND sg13g2_fill_1
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_13_989 VPWR VGND sg13g2_decap_8
XFILLER_32_1011 VPWR VGND sg13g2_decap_8
Xhold4 mac1.products_ff\[149\] VPWR VGND net44 sg13g2_dlygate4sd3_1
XFILLER_35_525 VPWR VGND sg13g2_decap_4
X_3990_ _0834_ _0788_ _0791_ _0831_ VPWR VGND sg13g2_and3_1
X_5660_ VGND VPWR _2369_ _2362_ _2359_ sg13g2_or2_1
X_4611_ _1426_ _1425_ _1422_ VPWR VGND sg13g2_nand2b_1
X_5591_ _2313_ _2311_ net28 VPWR VGND sg13g2_xor2_1
X_4542_ net830 net882 net833 _1360_ VPWR VGND net880 sg13g2_nand4_1
X_4473_ _1298_ _1293_ _1297_ VPWR VGND sg13g2_nand2_1
Xhold404 DP_2.matrix\[3\] VPWR VGND net444 sg13g2_dlygate4sd3_1
Xhold426 DP_2.matrix\[42\] VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold415 _2261_ VPWR VGND net455 sg13g2_dlygate4sd3_1
X_3424_ _0288_ net993 net927 VPWR VGND sg13g2_nand2_1
X_6212_ net1041 VGND VPWR net126 mac1.sum_lvl2_ff\[39\] clknet_leaf_62_clk sg13g2_dfrbpq_1
Xhold459 mac1.sum_lvl2_ff\[26\] VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold437 DP_1.matrix\[43\] VPWR VGND net477 sg13g2_dlygate4sd3_1
Xhold448 _2258_ VPWR VGND net488 sg13g2_dlygate4sd3_1
Xfanout906 net907 net906 VPWR VGND sg13g2_buf_8
X_6143_ net1061 VGND VPWR _0248_ DP_4.matrix\[4\] clknet_leaf_26_clk sg13g2_dfrbpq_1
Xfanout939 net940 net939 VPWR VGND sg13g2_buf_2
Xfanout917 DP_2.matrix\[38\] net917 VPWR VGND sg13g2_buf_1
X_3355_ _2941_ DP_2.matrix\[78\] net1007 VPWR VGND sg13g2_nand2_1
Xfanout928 net431 net928 VPWR VGND sg13g2_buf_8
X_3286_ _2875_ _2854_ _2874_ VPWR VGND sg13g2_xnor2_1
X_6074_ net1065 VGND VPWR _0202_ DP_2.matrix\[6\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_5025_ _1823_ _1817_ _1821_ VPWR VGND sg13g2_xnor2_1
X_5927_ net966 _0185_ VPWR VGND sg13g2_buf_1
X_5858_ net928 net757 _2551_ VPWR VGND sg13g2_nor2_1
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
X_5789_ net806 net779 _2495_ VPWR VGND sg13g2_nor2_1
X_4809_ _1619_ net877 DP_4.matrix\[6\] VPWR VGND sg13g2_nand2_2
XFILLER_49_628 VPWR VGND sg13g2_decap_8
XFILLER_45_867 VPWR VGND sg13g2_decap_8
XFILLER_44_344 VPWR VGND sg13g2_fill_2
XFILLER_44_95 VPWR VGND sg13g2_fill_1
XFILLER_44_73 VPWR VGND sg13g2_fill_2
XFILLER_8_278 VPWR VGND sg13g2_fill_2
XFILLER_5_930 VPWR VGND sg13g2_decap_8
X_3140_ _2721_ VPWR _2732_ VGND _2701_ _2722_ sg13g2_o21ai_1
X_3071_ _2665_ _2663_ _2664_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_878 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
X_5712_ net932 net776 _2420_ VPWR VGND sg13g2_nor2_1
X_3973_ _0774_ VPWR _0817_ VGND _0772_ _0775_ sg13g2_o21ai_1
X_5643_ mac1.total_sum\[14\] mac2.total_sum\[14\] _2355_ VPWR VGND sg13g2_nor2_1
X_5574_ _0053_ _2298_ net348 VPWR VGND sg13g2_xnor2_1
X_4525_ _1347_ _1341_ _1346_ VPWR VGND sg13g2_xnor2_1
Xhold201 mac2.sum_lvl2_ff\[52\] VPWR VGND net241 sg13g2_dlygate4sd3_1
Xhold223 mac2.products_ff\[12\] VPWR VGND net263 sg13g2_dlygate4sd3_1
Xhold212 mac2.products_ff\[138\] VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold234 DP_3.matrix\[77\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold256 DP_4.matrix\[76\] VPWR VGND net296 sg13g2_dlygate4sd3_1
X_4456_ _1281_ _1276_ _1279_ VPWR VGND sg13g2_xnor2_1
Xhold267 DP_2.matrix\[76\] VPWR VGND net307 sg13g2_dlygate4sd3_1
Xhold278 _2154_ VPWR VGND net318 sg13g2_dlygate4sd3_1
Xhold245 mac1.sum_lvl2_ff\[15\] VPWR VGND net285 sg13g2_dlygate4sd3_1
X_3407_ _2973_ VPWR _0272_ VGND _2971_ _2974_ sg13g2_o21ai_1
Xhold289 DP_3.matrix\[37\] VPWR VGND net329 sg13g2_dlygate4sd3_1
X_4387_ _1214_ _1207_ _1213_ VPWR VGND sg13g2_xnor2_1
X_3338_ _2923_ _2884_ _2925_ VPWR VGND sg13g2_xor2_1
X_6126_ net1054 VGND VPWR _0237_ DP_3.matrix\[73\] clknet_leaf_28_clk sg13g2_dfrbpq_1
Xfanout758 net759 net758 VPWR VGND sg13g2_buf_8
Xfanout769 _2447_ net769 VPWR VGND sg13g2_buf_8
X_6057_ net1040 VGND VPWR _0191_ DP_1.matrix\[75\] clknet_leaf_64_clk sg13g2_dfrbpq_2
X_3269_ VGND VPWR _2858_ _2857_ _2833_ sg13g2_or2_1
X_5008_ _1805_ _1804_ _1795_ _1807_ VPWR VGND sg13g2_a21o_1
XFILLER_39_694 VPWR VGND sg13g2_decap_4
XFILLER_14_539 VPWR VGND sg13g2_fill_1
XFILLER_26_377 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_10_701 VPWR VGND sg13g2_fill_2
XFILLER_2_922 VPWR VGND sg13g2_decap_8
XFILLER_1_465 VPWR VGND sg13g2_fill_1
XFILLER_2_999 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_17_300 VPWR VGND sg13g2_decap_4
XFILLER_41_892 VPWR VGND sg13g2_decap_8
XFILLER_9_565 VPWR VGND sg13g2_fill_1
X_5290_ _2079_ _2062_ _2080_ VPWR VGND sg13g2_xor2_1
X_4310_ _1139_ net811 net858 VPWR VGND sg13g2_nand2_1
X_4241_ _1070_ _1069_ _1060_ _1072_ VPWR VGND sg13g2_a21o_1
XFILLER_45_1021 VPWR VGND sg13g2_decap_8
X_4172_ _0989_ _1004_ _1005_ VPWR VGND sg13g2_nor2_1
X_3123_ _2713_ _2714_ _2708_ _2716_ VPWR VGND sg13g2_nand3_1
X_3054_ _2649_ _2642_ _2647_ _2648_ VPWR VGND sg13g2_and3_1
X_3956_ VGND VPWR _0800_ _0768_ _0766_ sg13g2_or2_1
XFILLER_32_892 VPWR VGND sg13g2_decap_8
X_3887_ _0729_ _0730_ _0732_ _0733_ VPWR VGND sg13g2_or3_1
X_5626_ _2339_ _2340_ _2341_ VPWR VGND sg13g2_nor2b_1
X_5557_ _0050_ net425 _2287_ VPWR VGND sg13g2_xnor2_1
X_4508_ _1331_ _1326_ _1329_ VPWR VGND sg13g2_xnor2_1
X_5488_ _2223_ _2227_ _2233_ _2234_ VPWR VGND sg13g2_nor3_1
X_4439_ VGND VPWR _1230_ _1232_ _1265_ _1264_ sg13g2_a21oi_1
XFILLER_47_918 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_fill_2
X_6109_ net1067 VGND VPWR net204 mac1.sum_lvl1_ff\[4\] clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_18_108 VPWR VGND sg13g2_fill_1
XFILLER_26_163 VPWR VGND sg13g2_fill_2
XFILLER_27_697 VPWR VGND sg13g2_fill_2
XFILLER_14_325 VPWR VGND sg13g2_fill_2
XFILLER_41_188 VPWR VGND sg13g2_decap_8
XFILLER_10_531 VPWR VGND sg13g2_fill_1
XFILLER_6_568 VPWR VGND sg13g2_fill_1
XFILLER_1_273 VPWR VGND sg13g2_fill_1
XFILLER_38_907 VPWR VGND sg13g2_decap_8
XFILLER_46_973 VPWR VGND sg13g2_decap_8
XFILLER_45_461 VPWR VGND sg13g2_fill_1
XFILLER_33_656 VPWR VGND sg13g2_fill_1
X_3810_ _0658_ net974 net915 VPWR VGND sg13g2_nand2_1
X_4790_ VGND VPWR _1562_ _1564_ _1601_ _1600_ sg13g2_a21oi_1
X_3741_ _0596_ _0591_ _0594_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_1020 VPWR VGND sg13g2_decap_8
X_3672_ _0529_ _0506_ _0530_ VPWR VGND sg13g2_nor2b_1
X_6460_ net1051 VGND VPWR net463 mac2.sum_lvl3_ff\[4\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5411_ _0017_ _2171_ net378 VPWR VGND sg13g2_xnor2_1
X_6391_ net1073 VGND VPWR net195 mac2.sum_lvl1_ff\[4\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5342_ _2119_ _2120_ _2121_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_5273_ _2063_ _2039_ _2064_ VPWR VGND sg13g2_xor2_1
X_4224_ _1055_ net870 net805 VPWR VGND sg13g2_nand2_1
X_4155_ _0989_ net363 net809 VPWR VGND sg13g2_nand2_1
X_3106_ _2696_ _2698_ _2699_ VPWR VGND sg13g2_nor2b_1
X_4086_ VGND VPWR _0867_ _0898_ _0927_ _0897_ sg13g2_a21oi_1
XFILLER_37_951 VPWR VGND sg13g2_decap_8
XFILLER_43_409 VPWR VGND sg13g2_fill_1
X_3037_ _2631_ _2630_ _2633_ VPWR VGND sg13g2_xor2_1
X_4988_ _1787_ _1785_ _1786_ VPWR VGND sg13g2_nand2b_1
X_3939_ _0781_ _0782_ _0763_ _0784_ VPWR VGND sg13g2_nand3_1
XFILLER_20_873 VPWR VGND sg13g2_fill_2
X_5609_ _2320_ _2323_ _2326_ _2328_ VPWR VGND sg13g2_or3_1
XFILLER_28_951 VPWR VGND sg13g2_decap_8
XFILLER_15_634 VPWR VGND sg13g2_fill_2
XFILLER_43_976 VPWR VGND sg13g2_decap_8
XFILLER_35_1020 VPWR VGND sg13g2_decap_8
Xinput16 uio_in[7] net16 VPWR VGND sg13g2_buf_1
XFILLER_7_811 VPWR VGND sg13g2_fill_2
XFILLER_11_895 VPWR VGND sg13g2_fill_2
XFILLER_37_236 VPWR VGND sg13g2_fill_1
XFILLER_38_759 VPWR VGND sg13g2_fill_1
X_5960_ net858 _0234_ VPWR VGND sg13g2_buf_1
XFILLER_19_973 VPWR VGND sg13g2_decap_8
XFILLER_46_781 VPWR VGND sg13g2_decap_4
X_5891_ net397 VPWR _0227_ VGND _2490_ _2572_ sg13g2_o21ai_1
X_4911_ net279 net800 _0089_ VPWR VGND sg13g2_and2_1
XFILLER_34_954 VPWR VGND sg13g2_decap_8
X_4842_ _1649_ _1640_ _1651_ VPWR VGND sg13g2_xor2_1
X_4773_ _1556_ VPWR _1584_ VGND _1550_ _1557_ sg13g2_o21ai_1
X_3724_ _0580_ _0552_ _0578_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_192 VPWR VGND sg13g2_fill_1
X_3655_ _0512_ _0509_ _0513_ VPWR VGND sg13g2_xor2_1
X_6443_ net1072 VGND VPWR net188 mac2.sum_lvl2_ff\[22\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_3586_ _0446_ DP_2.matrix\[3\] net982 VPWR VGND sg13g2_nand2_1
X_6374_ net1050 VGND VPWR _0092_ mac2.products_ff\[139\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5325_ _2100_ _2103_ _2106_ _2108_ VPWR VGND sg13g2_or3_1
X_5256_ _2046_ _2008_ _2048_ VPWR VGND sg13g2_xor2_1
X_4207_ _1028_ _1036_ _1038_ _1039_ VPWR VGND sg13g2_or3_1
X_5187_ VGND VPWR _1981_ _1980_ _1957_ sg13g2_or2_1
X_4138_ _0976_ net961 net1004 VPWR VGND sg13g2_nand2_1
X_4069_ _0885_ _0909_ _0910_ VPWR VGND sg13g2_nor2_1
XFILLER_28_269 VPWR VGND sg13g2_decap_8
XFILLER_12_604 VPWR VGND sg13g2_fill_1
XFILLER_19_1015 VPWR VGND sg13g2_decap_8
XFILLER_25_987 VPWR VGND sg13g2_decap_8
XFILLER_40_913 VPWR VGND sg13g2_decap_8
XFILLER_11_114 VPWR VGND sg13g2_fill_1
XFILLER_12_659 VPWR VGND sg13g2_decap_8
XFILLER_4_814 VPWR VGND sg13g2_decap_4
XFILLER_43_762 VPWR VGND sg13g2_fill_2
XFILLER_15_486 VPWR VGND sg13g2_decap_8
XFILLER_16_998 VPWR VGND sg13g2_decap_8
XFILLER_31_913 VPWR VGND sg13g2_decap_8
X_3440_ _0293_ _0301_ _0303_ _0304_ VPWR VGND sg13g2_or3_1
X_3371_ _2956_ net943 net1003 VPWR VGND sg13g2_nand2_1
X_6090_ net1040 VGND VPWR _0213_ DP_2.matrix\[73\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_5110_ _1906_ net848 net783 VPWR VGND sg13g2_nand2_1
X_5041_ _1836_ _1837_ _1831_ _1839_ VPWR VGND sg13g2_nand3_1
XFILLER_26_2 VPWR VGND sg13g2_fill_1
X_5943_ net910 _0209_ VPWR VGND sg13g2_buf_1
XFILLER_22_913 VPWR VGND sg13g2_decap_4
X_5874_ _2470_ _2468_ _2561_ VPWR VGND sg13g2_xor2_1
XFILLER_40_209 VPWR VGND sg13g2_fill_1
X_4825_ _0140_ _1633_ _1634_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_990 VPWR VGND sg13g2_decap_8
X_4756_ _1568_ _1522_ _1525_ _1565_ VPWR VGND sg13g2_and3_1
X_3707_ VGND VPWR _0503_ _0562_ _0564_ _0563_ sg13g2_a21oi_1
X_4687_ net825 net879 net823 net877 _1500_ VPWR VGND sg13g2_and4_1
X_3638_ _0495_ _0472_ _0497_ VPWR VGND sg13g2_xor2_1
X_6426_ net1059 VGND VPWR net133 mac2.sum_lvl2_ff\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_3569_ _0114_ _0384_ _0428_ VPWR VGND sg13g2_xnor2_1
X_6357_ net1059 VGND VPWR _0081_ mac2.products_ff\[70\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5308_ _2092_ VPWR _2094_ VGND _2091_ _2093_ sg13g2_o21ai_1
X_6288_ net1051 VGND VPWR net158 mac1.sum_lvl3_ff\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5239_ _1974_ _2031_ _2032_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_567 VPWR VGND sg13g2_fill_1
XFILLER_13_924 VPWR VGND sg13g2_fill_1
XFILLER_9_917 VPWR VGND sg13g2_fill_1
XFILLER_13_968 VPWR VGND sg13g2_decap_8
XFILLER_40_776 VPWR VGND sg13g2_fill_1
XFILLER_8_449 VPWR VGND sg13g2_fill_1
XFILLER_21_990 VPWR VGND sg13g2_decap_8
XFILLER_40_798 VPWR VGND sg13g2_fill_2
Xhold5 mac2.products_ff\[1\] VPWR VGND net45 sg13g2_dlygate4sd3_1
XFILLER_48_898 VPWR VGND sg13g2_decap_8
X_4610_ _1424_ _1391_ _1425_ VPWR VGND sg13g2_xor2_1
X_5590_ _2313_ mac1.total_sum\[3\] mac2.total_sum\[3\] VPWR VGND sg13g2_xnor2_1
X_4541_ net833 net829 net882 net880 _1359_ VPWR VGND sg13g2_and4_1
Xhold427 DP_4.matrix\[42\] VPWR VGND net467 sg13g2_dlygate4sd3_1
XFILLER_8_994 VPWR VGND sg13g2_decap_8
Xhold416 _0058_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold405 DP_1.matrix\[8\] VPWR VGND net445 sg13g2_dlygate4sd3_1
X_4472_ VGND VPWR _1296_ _1297_ _1295_ _1237_ sg13g2_a21oi_2
X_3423_ _0279_ VPWR _0287_ VGND _0271_ _0281_ sg13g2_o21ai_1
X_6211_ net1041 VGND VPWR net148 mac1.sum_lvl2_ff\[38\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xhold449 _0057_ VPWR VGND net489 sg13g2_dlygate4sd3_1
Xhold438 mac1.sum_lvl2_ff\[13\] VPWR VGND net478 sg13g2_dlygate4sd3_1
Xfanout907 net464 net907 VPWR VGND sg13g2_buf_8
X_6142_ net1096 VGND VPWR net80 mac1.sum_lvl1_ff\[15\] clknet_leaf_40_clk sg13g2_dfrbpq_1
Xfanout918 net442 net918 VPWR VGND sg13g2_buf_8
Xfanout929 net444 net929 VPWR VGND sg13g2_buf_8
X_3354_ _2940_ net888 net1007 VPWR VGND sg13g2_nand2_1
X_6073_ net1015 VGND VPWR _0103_ mac1.products_ff\[144\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3285_ _2872_ _2861_ _2874_ VPWR VGND sg13g2_xor2_1
X_5024_ _1817_ _1821_ _1822_ VPWR VGND sg13g2_and2_1
X_5926_ net968 _0184_ VPWR VGND sg13g2_buf_1
XFILLER_22_754 VPWR VGND sg13g2_fill_2
X_5857_ VGND VPWR net753 _2550_ _0199_ _2549_ sg13g2_a21oi_1
X_5788_ _2494_ net786 net766 VPWR VGND sg13g2_nand2_1
X_4808_ _1618_ net881 net996 VPWR VGND sg13g2_nand2_1
XFILLER_5_408 VPWR VGND sg13g2_fill_2
X_4739_ _1508_ VPWR _1551_ VGND _1506_ _1509_ sg13g2_o21ai_1
X_6409_ net1071 VGND VPWR net218 mac2.sum_lvl1_ff\[42\] clknet_leaf_41_clk sg13g2_dfrbpq_1
XFILLER_49_607 VPWR VGND sg13g2_decap_8
XFILLER_0_113 VPWR VGND sg13g2_fill_1
XFILLER_13_710 VPWR VGND sg13g2_fill_2
XFILLER_44_63 VPWR VGND sg13g2_fill_2
XFILLER_40_584 VPWR VGND sg13g2_decap_8
XFILLER_5_986 VPWR VGND sg13g2_decap_8
X_3070_ _2664_ net958 net889 VPWR VGND sg13g2_nand2_2
XFILLER_48_684 VPWR VGND sg13g2_fill_1
XFILLER_35_312 VPWR VGND sg13g2_fill_2
XFILLER_39_1007 VPWR VGND sg13g2_decap_8
XFILLER_23_529 VPWR VGND sg13g2_decap_8
X_5711_ _2419_ net770 _2418_ net763 net277 VPWR VGND sg13g2_a22oi_1
X_3972_ _0816_ _0811_ _0815_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_551 VPWR VGND sg13g2_fill_1
X_5642_ _2354_ mac1.total_sum\[14\] mac2.total_sum\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_31_584 VPWR VGND sg13g2_decap_4
X_5573_ net347 mac2.sum_lvl3_ff\[34\] _2301_ VPWR VGND sg13g2_xor2_1
X_4524_ _1346_ _1333_ _1345_ VPWR VGND sg13g2_xnor2_1
Xhold202 mac1.sum_lvl1_ff\[49\] VPWR VGND net242 sg13g2_dlygate4sd3_1
Xhold224 mac2.products_ff\[15\] VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold235 DP_2.matrix\[80\] VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold213 mac2.products_ff\[0\] VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold268 DP_3.matrix\[78\] VPWR VGND net308 sg13g2_dlygate4sd3_1
X_4455_ _1280_ _1279_ _1276_ VPWR VGND sg13g2_nand2b_1
Xhold257 DP_1.matrix\[76\] VPWR VGND net297 sg13g2_dlygate4sd3_1
Xhold246 _2138_ VPWR VGND net286 sg13g2_dlygate4sd3_1
Xhold279 _0027_ VPWR VGND net319 sg13g2_dlygate4sd3_1
X_3406_ VGND VPWR _0271_ _0270_ _0268_ sg13g2_or2_1
X_4386_ _1212_ _1208_ _1213_ VPWR VGND sg13g2_xor2_1
X_3337_ _2884_ _2923_ _2924_ VPWR VGND sg13g2_nor2_1
X_6125_ net1054 VGND VPWR _0236_ DP_3.matrix\[72\] clknet_leaf_15_clk sg13g2_dfrbpq_2
Xfanout759 net762 net759 VPWR VGND sg13g2_buf_8
X_6056_ net1041 VGND VPWR _0190_ DP_1.matrix\[74\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_3268_ _2857_ net895 net1006 VPWR VGND sg13g2_nand2_1
XFILLER_22_1011 VPWR VGND sg13g2_decap_8
XFILLER_27_802 VPWR VGND sg13g2_fill_1
XFILLER_39_662 VPWR VGND sg13g2_fill_1
X_3199_ _2759_ VPWR _2790_ VGND _2750_ _2760_ sg13g2_o21ai_1
XFILLER_38_172 VPWR VGND sg13g2_fill_2
X_5007_ _1804_ _1805_ _1795_ _1806_ VPWR VGND sg13g2_nand3_1
XFILLER_27_868 VPWR VGND sg13g2_decap_8
X_5909_ _2584_ net821 net760 VPWR VGND sg13g2_nand2_1
XFILLER_30_43 VPWR VGND sg13g2_fill_1
XFILLER_2_978 VPWR VGND sg13g2_decap_8
XFILLER_39_30 VPWR VGND sg13g2_fill_2
XFILLER_49_437 VPWR VGND sg13g2_fill_1
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_312 VPWR VGND sg13g2_fill_1
XFILLER_41_871 VPWR VGND sg13g2_decap_8
XFILLER_9_511 VPWR VGND sg13g2_fill_1
XFILLER_45_1000 VPWR VGND sg13g2_decap_8
X_4240_ _1069_ _1070_ _1060_ _1071_ VPWR VGND sg13g2_nand3_1
X_4171_ _1004_ net870 net808 VPWR VGND sg13g2_nand2_2
X_3122_ _2715_ _2708_ _2713_ _2714_ VPWR VGND sg13g2_and3_1
XFILLER_49_982 VPWR VGND sg13g2_decap_8
X_3053_ _2643_ VPWR _2648_ VGND _2644_ _2646_ sg13g2_o21ai_1
XFILLER_35_131 VPWR VGND sg13g2_fill_2
X_3955_ _0758_ VPWR _0799_ VGND _0717_ _0756_ sg13g2_o21ai_1
XFILLER_32_871 VPWR VGND sg13g2_decap_8
X_3886_ _0732_ net960 net922 net963 net919 VPWR VGND sg13g2_a22oi_1
X_5625_ VGND VPWR _2340_ mac2.total_sum\[11\] mac1.total_sum\[11\] sg13g2_or2_1
X_5556_ VGND VPWR net381 _2283_ _2287_ _2280_ sg13g2_a21oi_1
X_4507_ _1330_ _1329_ _1326_ VPWR VGND sg13g2_nand2b_1
X_5487_ _2233_ _2226_ _2231_ VPWR VGND sg13g2_nand2_1
X_4438_ _1262_ _1240_ _1264_ VPWR VGND sg13g2_xor2_1
X_4369_ _1197_ _1164_ _1196_ VPWR VGND sg13g2_nand2b_1
X_6108_ net1061 VGND VPWR _0225_ DP_3.matrix\[5\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_6039_ net1047 VGND VPWR _0176_ DP_1.matrix\[4\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_27_632 VPWR VGND sg13g2_fill_2
XFILLER_25_65 VPWR VGND sg13g2_fill_2
XFILLER_10_565 VPWR VGND sg13g2_fill_2
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_952 VPWR VGND sg13g2_decap_8
XFILLER_18_643 VPWR VGND sg13g2_fill_1
XFILLER_45_484 VPWR VGND sg13g2_fill_2
XFILLER_18_698 VPWR VGND sg13g2_fill_2
XFILLER_33_624 VPWR VGND sg13g2_decap_4
X_3740_ _0595_ _0594_ _0591_ VPWR VGND sg13g2_nand2b_1
XFILLER_32_189 VPWR VGND sg13g2_decap_4
XFILLER_9_363 VPWR VGND sg13g2_fill_1
X_3671_ _0529_ _0507_ _0528_ VPWR VGND sg13g2_xnor2_1
X_5410_ _2174_ _2171_ _2173_ VPWR VGND sg13g2_nand2b_1
X_6390_ net1072 VGND VPWR net78 mac2.sum_lvl1_ff\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5341_ VGND VPWR _2120_ mac1.sum_lvl2_ff\[11\] mac1.sum_lvl2_ff\[30\] sg13g2_or2_1
X_5272_ _2063_ net783 net997 VPWR VGND sg13g2_nand2_1
X_4223_ _1037_ VPWR _1054_ VGND _1028_ _1038_ sg13g2_o21ai_1
X_4154_ _0987_ _0981_ _0081_ VPWR VGND sg13g2_xor2_1
X_3105_ VGND VPWR _2698_ _2697_ _2664_ sg13g2_or2_1
X_4085_ _0924_ _0923_ _0926_ VPWR VGND sg13g2_xor2_1
X_3036_ _2632_ _2630_ _2631_ VPWR VGND sg13g2_nand2_1
XFILLER_37_930 VPWR VGND sg13g2_decap_8
XFILLER_36_451 VPWR VGND sg13g2_fill_1
XFILLER_36_473 VPWR VGND sg13g2_fill_1
XFILLER_24_668 VPWR VGND sg13g2_fill_2
X_4987_ _1786_ net854 net783 VPWR VGND sg13g2_nand2_1
X_3938_ _0783_ _0763_ _0781_ _0782_ VPWR VGND sg13g2_and3_1
X_3869_ _0692_ VPWR _0715_ VGND _0657_ _0690_ sg13g2_o21ai_1
X_5608_ _2326_ VPWR _2327_ VGND _2320_ _2323_ sg13g2_o21ai_1
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
X_5539_ _2272_ net540 _0061_ VPWR VGND sg13g2_and2_1
XFILLER_28_930 VPWR VGND sg13g2_decap_8
XFILLER_43_955 VPWR VGND sg13g2_decap_8
XFILLER_7_834 VPWR VGND sg13g2_fill_2
XFILLER_19_930 VPWR VGND sg13g2_fill_1
XFILLER_38_749 VPWR VGND sg13g2_fill_2
X_4910_ _0144_ _1708_ _1715_ VPWR VGND sg13g2_xnor2_1
X_5890_ _2483_ _2485_ _2572_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_933 VPWR VGND sg13g2_decap_8
X_4841_ _1649_ _1640_ _1650_ VPWR VGND sg13g2_nor2b_1
X_4772_ _1581_ _1573_ _1583_ VPWR VGND sg13g2_xor2_1
X_3723_ _0579_ _0578_ _0552_ VPWR VGND sg13g2_nand2b_1
X_3654_ _0512_ _0487_ _0510_ VPWR VGND sg13g2_xnor2_1
X_6442_ net1059 VGND VPWR net155 mac2.sum_lvl2_ff\[21\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_3585_ _0445_ DP_2.matrix\[4\] net982 VPWR VGND sg13g2_nand2_1
X_6373_ net1050 VGND VPWR _0091_ mac2.products_ff\[138\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5324_ _2106_ VPWR _2107_ VGND _2100_ _2103_ sg13g2_o21ai_1
X_5255_ _2008_ _2046_ _2047_ VPWR VGND sg13g2_nor2_1
X_4206_ VGND VPWR _1034_ _1035_ _1038_ _1029_ sg13g2_a21oi_1
X_5186_ _1980_ net789 net997 VPWR VGND sg13g2_nand2_1
XFILLER_29_705 VPWR VGND sg13g2_fill_2
XFILLER_29_738 VPWR VGND sg13g2_fill_2
X_4137_ _0963_ VPWR _0975_ VGND _0936_ _0961_ sg13g2_o21ai_1
XFILLER_29_749 VPWR VGND sg13g2_fill_2
X_4068_ _0909_ net964 net906 VPWR VGND sg13g2_nand2_2
X_3019_ _0067_ _2601_ _2614_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_966 VPWR VGND sg13g2_decap_8
XFILLER_40_969 VPWR VGND sg13g2_decap_8
XFILLER_47_74 VPWR VGND sg13g2_fill_2
XFILLER_15_432 VPWR VGND sg13g2_fill_1
XFILLER_16_977 VPWR VGND sg13g2_decap_8
XFILLER_31_969 VPWR VGND sg13g2_decap_8
XFILLER_6_152 VPWR VGND sg13g2_fill_1
XFILLER_6_141 VPWR VGND sg13g2_fill_1
X_3370_ _2943_ VPWR _2955_ VGND _2917_ _2940_ sg13g2_o21ai_1
X_5040_ _1838_ _1831_ _1836_ _1837_ VPWR VGND sg13g2_and3_1
XFILLER_38_502 VPWR VGND sg13g2_decap_4
XFILLER_38_546 VPWR VGND sg13g2_decap_4
XFILLER_38_579 VPWR VGND sg13g2_fill_2
X_5942_ net912 _0208_ VPWR VGND sg13g2_buf_1
X_5873_ _2560_ VPWR _0221_ VGND net758 _2559_ sg13g2_o21ai_1
XFILLER_22_969 VPWR VGND sg13g2_decap_8
X_4824_ VGND VPWR _1603_ _1606_ _1634_ _1601_ sg13g2_a21oi_1
X_4755_ _1525_ _1522_ _1565_ _1567_ VPWR VGND sg13g2_a21o_1
X_3706_ _0533_ VPWR _0563_ VGND _0501_ _0532_ sg13g2_o21ai_1
X_4686_ _1499_ net823 net877 VPWR VGND sg13g2_nand2_1
X_3637_ _0496_ _0472_ _0495_ VPWR VGND sg13g2_nand2_1
X_6425_ net1058 VGND VPWR net244 mac2.sum_lvl2_ff\[1\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_1_807 VPWR VGND sg13g2_fill_1
X_3568_ _0383_ _0428_ _0382_ _0429_ VPWR VGND sg13g2_nand3_1
X_6356_ net1052 VGND VPWR _0080_ mac2.products_ff\[69\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5307_ net495 _2091_ _0009_ VPWR VGND sg13g2_xor2_1
X_3499_ _0329_ VPWR _0361_ VGND _0327_ _0330_ sg13g2_o21ai_1
X_6287_ net1025 VGND VPWR net55 mac1.sum_lvl3_ff\[32\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5238_ VGND VPWR _1970_ _2003_ _2031_ _2002_ sg13g2_a21oi_1
X_5169_ _1962_ _1954_ _1964_ VPWR VGND sg13g2_xor2_1
XFILLER_44_505 VPWR VGND sg13g2_fill_2
XFILLER_17_99 VPWR VGND sg13g2_fill_2
XFILLER_24_262 VPWR VGND sg13g2_fill_2
XFILLER_13_947 VPWR VGND sg13g2_decap_8
XFILLER_3_188 VPWR VGND sg13g2_decap_8
Xhold6 mac1.sum_lvl1_ff\[46\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_877 VPWR VGND sg13g2_decap_8
XFILLER_43_582 VPWR VGND sg13g2_decap_4
XFILLER_30_232 VPWR VGND sg13g2_fill_1
XFILLER_31_788 VPWR VGND sg13g2_fill_1
XFILLER_8_973 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_4_3_0_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_4540_ _1358_ net884 net827 VPWR VGND sg13g2_nand2_1
Xhold406 _0160_ VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold417 mac2.sum_lvl3_ff\[6\] VPWR VGND net457 sg13g2_dlygate4sd3_1
X_4471_ _1266_ VPWR _1296_ VGND _1235_ _1265_ sg13g2_o21ai_1
X_3422_ _0285_ _2982_ _0073_ VPWR VGND sg13g2_xor2_1
Xhold439 _2130_ VPWR VGND net479 sg13g2_dlygate4sd3_1
Xhold428 mac1.sum_lvl2_ff\[14\] VPWR VGND net468 sg13g2_dlygate4sd3_1
X_6210_ net1084 VGND VPWR net215 mac1.sum_lvl2_ff\[34\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6141_ net1061 VGND VPWR net351 DP_4.matrix\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_2
Xfanout919 net920 net919 VPWR VGND sg13g2_buf_2
X_3353_ _2939_ net945 net1003 VPWR VGND sg13g2_nand2_1
Xfanout908 net909 net908 VPWR VGND sg13g2_buf_8
X_3284_ _2861_ _2872_ _2873_ VPWR VGND sg13g2_nor2_1
X_6072_ net1065 VGND VPWR _0201_ DP_2.matrix\[5\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_5023_ _1818_ _1820_ _1821_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_888 VPWR VGND sg13g2_decap_8
XFILLER_0_1011 VPWR VGND sg13g2_decap_8
XFILLER_19_590 VPWR VGND sg13g2_decap_8
X_5925_ net971 _0183_ VPWR VGND sg13g2_buf_1
X_5856_ _2429_ _2417_ _2550_ VPWR VGND sg13g2_xor2_1
X_4807_ VGND VPWR _1617_ _1590_ _1588_ sg13g2_or2_1
XFILLER_16_1019 VPWR VGND sg13g2_decap_8
X_5787_ VGND VPWR _2593_ net777 _2493_ _2492_ sg13g2_a21oi_1
X_2999_ net903 net956 net898 net954 _2597_ VPWR VGND sg13g2_and4_1
X_4738_ _1550_ _1545_ _1549_ VPWR VGND sg13g2_xnor2_1
X_4669_ _1482_ _1419_ _1483_ VPWR VGND sg13g2_xor2_1
X_6408_ net1073 VGND VPWR net229 mac2.sum_lvl1_ff\[41\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_6339_ net1055 VGND VPWR _0084_ mac2.products_ff\[0\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_28_32 VPWR VGND sg13g2_fill_1
XFILLER_44_346 VPWR VGND sg13g2_fill_1
XFILLER_44_75 VPWR VGND sg13g2_fill_1
XFILLER_13_799 VPWR VGND sg13g2_fill_2
XFILLER_5_910 VPWR VGND sg13g2_fill_1
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_4_497 VPWR VGND sg13g2_fill_2
XFILLER_39_129 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_59_clk clknet_4_9_0_clk clknet_leaf_59_clk VPWR VGND sg13g2_buf_8
X_3971_ _0815_ _0765_ _0812_ VPWR VGND sg13g2_xnor2_1
X_5710_ net924 net937 net774 _2418_ VPWR VGND sg13g2_mux2_1
X_5641_ VGND VPWR mac1.total_sum\[13\] mac2.total_sum\[13\] _2353_ _2351_ sg13g2_a21oi_1
X_5572_ mac2.sum_lvl3_ff\[34\] net347 _2300_ VPWR VGND sg13g2_nor2_1
X_4523_ _1345_ _1342_ _1344_ VPWR VGND sg13g2_xnor2_1
Xhold225 mac1.sum_lvl2_ff\[0\] VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold214 mac2.products_ff\[6\] VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold203 mac2.sum_lvl1_ff\[85\] VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold269 DP_4.matrix\[79\] VPWR VGND net309 sg13g2_dlygate4sd3_1
Xhold258 DP_3.matrix\[79\] VPWR VGND net298 sg13g2_dlygate4sd3_1
X_4454_ _1278_ _1252_ _1279_ VPWR VGND sg13g2_xor2_1
Xhold236 DP_1.matrix\[74\] VPWR VGND net276 sg13g2_dlygate4sd3_1
Xhold247 _0006_ VPWR VGND net287 sg13g2_dlygate4sd3_1
X_3405_ _2969_ _0269_ _0270_ VPWR VGND sg13g2_nor2_1
X_4385_ _1212_ _1169_ _1210_ VPWR VGND sg13g2_xnor2_1
X_3336_ _2923_ _2914_ _2922_ VPWR VGND sg13g2_xnor2_1
X_6124_ net1070 VGND VPWR net65 mac1.sum_lvl1_ff\[9\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_6055_ net1023 VGND VPWR _0066_ mac1.products_ff\[138\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_3267_ _2856_ net890 net945 VPWR VGND sg13g2_nand2_1
X_5006_ _1802_ _1801_ _1796_ _1805_ VPWR VGND sg13g2_a21o_1
X_3198_ _2787_ _2779_ _2789_ VPWR VGND sg13g2_xor2_1
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_35_880 VPWR VGND sg13g2_decap_8
XFILLER_41_349 VPWR VGND sg13g2_fill_2
X_5908_ _2520_ _2516_ _2583_ VPWR VGND sg13g2_xor2_1
X_5839_ _2400_ _2378_ _2539_ VPWR VGND sg13g2_xor2_1
XFILLER_5_239 VPWR VGND sg13g2_fill_2
XFILLER_2_957 VPWR VGND sg13g2_decap_8
XFILLER_7_1006 VPWR VGND sg13g2_decap_8
XFILLER_39_42 VPWR VGND sg13g2_fill_1
XFILLER_17_357 VPWR VGND sg13g2_decap_4
XFILLER_26_880 VPWR VGND sg13g2_decap_8
X_4170_ _1003_ net808 DP_3.matrix\[36\] net809 net870 VPWR VGND sg13g2_a22oi_1
X_3121_ _2709_ VPWR _2714_ VGND _2710_ _2712_ sg13g2_o21ai_1
XFILLER_1_990 VPWR VGND sg13g2_decap_8
XFILLER_49_961 VPWR VGND sg13g2_decap_8
X_3052_ _2643_ _2644_ _2646_ _2647_ VPWR VGND sg13g2_or3_1
XFILLER_35_121 VPWR VGND sg13g2_fill_2
X_3954_ _0784_ VPWR _0798_ VGND _0762_ _0785_ sg13g2_o21ai_1
XFILLER_23_349 VPWR VGND sg13g2_fill_1
X_3885_ net919 net963 net922 _0731_ VPWR VGND net960 sg13g2_nand4_1
X_5624_ mac1.total_sum\[11\] mac2.total_sum\[11\] _2339_ VPWR VGND sg13g2_and2_1
X_5555_ net424 _2285_ _2286_ VPWR VGND sg13g2_nor2b_1
X_4506_ _1328_ _1303_ _1329_ VPWR VGND sg13g2_xor2_1
XFILLER_2_209 VPWR VGND sg13g2_fill_2
X_5486_ _0034_ _2231_ _2232_ VPWR VGND sg13g2_xnor2_1
X_4437_ _1262_ _1240_ _1263_ VPWR VGND sg13g2_nor2b_1
X_6107_ net1061 VGND VPWR _0224_ DP_3.matrix\[4\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_4368_ _1196_ _1165_ _1194_ VPWR VGND sg13g2_xnor2_1
X_3319_ VGND VPWR _2847_ _2879_ _2907_ _2878_ sg13g2_a21oi_1
X_4299_ _1128_ _1120_ _1126_ VPWR VGND sg13g2_xnor2_1
X_6038_ net1044 VGND VPWR _0175_ DP_1.matrix\[3\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_14_327 VPWR VGND sg13g2_fill_1
XFILLER_10_588 VPWR VGND sg13g2_fill_2
XFILLER_41_87 VPWR VGND sg13g2_decap_8
XFILLER_29_1007 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_fill_2
XFILLER_18_611 VPWR VGND sg13g2_decap_8
XFILLER_46_931 VPWR VGND sg13g2_decap_8
XFILLER_18_666 VPWR VGND sg13g2_fill_1
XFILLER_32_102 VPWR VGND sg13g2_fill_2
XFILLER_20_319 VPWR VGND sg13g2_fill_1
X_3670_ _0526_ _0514_ _0528_ VPWR VGND sg13g2_xor2_1
X_5340_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] _2119_ VPWR VGND sg13g2_and2_1
X_5271_ _2062_ net782 net997 VPWR VGND sg13g2_nand2_1
X_4222_ _1051_ _1050_ _1053_ VPWR VGND sg13g2_xor2_1
XFILLER_29_909 VPWR VGND sg13g2_decap_8
X_4153_ _0988_ _0981_ _0987_ VPWR VGND sg13g2_nand2_1
X_3104_ _2697_ net957 net887 VPWR VGND sg13g2_nand2_1
X_4084_ VGND VPWR _0925_ _0924_ _0923_ sg13g2_or2_1
X_3035_ _2631_ _2611_ _2613_ VPWR VGND sg13g2_nand2_1
XFILLER_36_463 VPWR VGND sg13g2_fill_1
XFILLER_37_986 VPWR VGND sg13g2_decap_8
XFILLER_23_146 VPWR VGND sg13g2_fill_2
X_4986_ _1762_ VPWR _1785_ VGND _1739_ _1760_ sg13g2_o21ai_1
X_3937_ _0770_ VPWR _0782_ VGND _0778_ _0780_ sg13g2_o21ai_1
X_3868_ _0706_ VPWR _0714_ VGND _0686_ _0707_ sg13g2_o21ai_1
XFILLER_20_875 VPWR VGND sg13g2_fill_1
X_3799_ _0646_ _0645_ _0640_ _0648_ VPWR VGND sg13g2_a21o_1
X_5607_ mac2.total_sum\[7\] mac1.total_sum\[7\] _2326_ VPWR VGND sg13g2_xor2_1
X_5538_ _2265_ _2268_ _2271_ _2273_ VPWR VGND sg13g2_or3_1
X_5469_ _2219_ mac2.sum_lvl2_ff\[27\] mac2.sum_lvl2_ff\[8\] VPWR VGND sg13g2_xnor2_1
XFILLER_47_706 VPWR VGND sg13g2_fill_2
XFILLER_27_452 VPWR VGND sg13g2_decap_4
XFILLER_28_986 VPWR VGND sg13g2_decap_8
XFILLER_43_934 VPWR VGND sg13g2_decap_8
XFILLER_42_422 VPWR VGND sg13g2_fill_2
XFILLER_42_444 VPWR VGND sg13g2_fill_2
XFILLER_11_875 VPWR VGND sg13g2_fill_2
XFILLER_6_367 VPWR VGND sg13g2_fill_2
XFILLER_42_1015 VPWR VGND sg13g2_decap_8
XFILLER_38_739 VPWR VGND sg13g2_fill_1
XFILLER_46_772 VPWR VGND sg13g2_fill_1
XFILLER_34_912 VPWR VGND sg13g2_decap_8
X_4840_ _1649_ _1641_ _1648_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_606 VPWR VGND sg13g2_fill_1
XFILLER_21_628 VPWR VGND sg13g2_decap_8
XFILLER_33_466 VPWR VGND sg13g2_fill_2
XFILLER_34_989 VPWR VGND sg13g2_decap_8
X_4771_ _1581_ _1573_ _1582_ VPWR VGND sg13g2_nor2b_1
X_3722_ _0576_ _0538_ _0578_ VPWR VGND sg13g2_xor2_1
X_3653_ VGND VPWR _0511_ _0510_ _0487_ sg13g2_or2_1
X_6441_ net1058 VGND VPWR net119 mac2.sum_lvl2_ff\[20\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6372_ net1050 VGND VPWR net290 mac2.products_ff\[137\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5323_ mac1.sum_lvl2_ff\[7\] mac1.sum_lvl2_ff\[26\] _2106_ VPWR VGND sg13g2_xor2_1
X_3584_ _0444_ net986 net927 VPWR VGND sg13g2_nand2_1
X_5254_ _2046_ _2037_ _2045_ VPWR VGND sg13g2_xnor2_1
X_5185_ _1979_ net785 net841 VPWR VGND sg13g2_nand2_1
X_4205_ _1034_ _1035_ _1029_ _1037_ VPWR VGND sg13g2_nand3_1
X_4136_ VGND VPWR _0944_ _0967_ _0974_ _0969_ sg13g2_a21oi_1
X_4067_ _0908_ net968 net1004 VPWR VGND sg13g2_nand2_1
X_3018_ _2601_ _2614_ _2615_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_934 VPWR VGND sg13g2_decap_8
X_4969_ _1765_ _1766_ _1768_ _1769_ VPWR VGND sg13g2_or3_1
XFILLER_40_948 VPWR VGND sg13g2_decap_8
XFILLER_47_536 VPWR VGND sg13g2_fill_2
XFILLER_43_720 VPWR VGND sg13g2_fill_2
XFILLER_16_956 VPWR VGND sg13g2_decap_8
XFILLER_43_764 VPWR VGND sg13g2_fill_1
XFILLER_31_948 VPWR VGND sg13g2_decap_8
XFILLER_6_175 VPWR VGND sg13g2_fill_2
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
X_5941_ net914 _0207_ VPWR VGND sg13g2_buf_1
XFILLER_46_580 VPWR VGND sg13g2_fill_2
X_5872_ _2560_ net884 net758 VPWR VGND sg13g2_nand2_1
XFILLER_21_436 VPWR VGND sg13g2_fill_2
X_4823_ _1631_ _1632_ _1633_ VPWR VGND sg13g2_nor2b_1
X_4754_ VGND VPWR _1522_ _1525_ _1566_ _1565_ sg13g2_a21oi_1
X_3705_ _0504_ _0561_ _0562_ VPWR VGND sg13g2_nor2b_1
X_4685_ _1498_ net881 net822 VPWR VGND sg13g2_nand2_1
X_3636_ _0494_ _0483_ _0495_ VPWR VGND sg13g2_xor2_1
X_6424_ net1057 VGND VPWR net47 mac2.sum_lvl2_ff\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_3567_ _0426_ _0427_ _0428_ VPWR VGND sg13g2_and2_1
X_6355_ net1051 VGND VPWR _0079_ mac2.products_ff\[68\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5306_ _2093_ mac1.sum_lvl2_ff\[22\] net494 VPWR VGND sg13g2_xnor2_1
X_6286_ net1024 VGND VPWR net53 mac1.sum_lvl3_ff\[31\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_5237_ _2028_ _2027_ _2030_ VPWR VGND sg13g2_xor2_1
XFILLER_0_329 VPWR VGND sg13g2_fill_2
X_3498_ _0360_ _0355_ _0359_ VPWR VGND sg13g2_xnor2_1
X_5168_ _1963_ _1954_ _1962_ VPWR VGND sg13g2_nand2b_1
X_4119_ _0942_ _0934_ _0941_ _0958_ VPWR VGND sg13g2_a21o_1
X_5099_ _1894_ _1895_ _1893_ _1896_ VPWR VGND sg13g2_nand3_1
XFILLER_44_517 VPWR VGND sg13g2_fill_1
XFILLER_32_1025 VPWR VGND sg13g2_decap_4
XFILLER_48_812 VPWR VGND sg13g2_fill_1
XFILLER_0_885 VPWR VGND sg13g2_decap_8
Xhold7 mac2.sum_lvl1_ff\[0\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_48_856 VPWR VGND sg13g2_decap_8
XFILLER_47_355 VPWR VGND sg13g2_fill_2
XFILLER_12_992 VPWR VGND sg13g2_decap_8
XFILLER_8_952 VPWR VGND sg13g2_decap_8
Xhold407 DP_3.matrix\[43\] VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold418 _2266_ VPWR VGND net458 sg13g2_dlygate4sd3_1
X_4470_ _1238_ _1294_ _1295_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_1010 VPWR VGND sg13g2_decap_8
X_3421_ _2982_ _0285_ _0286_ VPWR VGND sg13g2_and2_1
Xhold429 _2136_ VPWR VGND net469 sg13g2_dlygate4sd3_1
X_3352_ _2922_ _2914_ _2921_ _2938_ VPWR VGND sg13g2_a21o_1
X_6140_ net1060 VGND VPWR _0246_ DP_4.matrix\[2\] clknet_leaf_27_clk sg13g2_dfrbpq_1
Xfanout909 net466 net909 VPWR VGND sg13g2_buf_8
X_3283_ _2870_ _2862_ _2872_ VPWR VGND sg13g2_xor2_1
X_6071_ net1047 VGND VPWR _0200_ DP_2.matrix\[4\] clknet_leaf_57_clk sg13g2_dfrbpq_2
X_5022_ VGND VPWR _1820_ _1819_ _1786_ sg13g2_or2_1
XFILLER_38_311 VPWR VGND sg13g2_fill_1
XFILLER_17_0 VPWR VGND sg13g2_fill_1
XFILLER_39_867 VPWR VGND sg13g2_decap_8
X_5924_ net974 _0182_ VPWR VGND sg13g2_buf_1
X_5855_ net929 net753 _2549_ VPWR VGND sg13g2_nor2_1
X_4806_ _1578_ VPWR _1616_ VGND _1575_ _1579_ sg13g2_o21ai_1
X_5786_ net768 VPWR _2492_ VGND net996 net777 sg13g2_o21ai_1
X_2998_ net958 net896 _2596_ VPWR VGND sg13g2_and2_1
X_4737_ _1549_ _1499_ _1546_ VPWR VGND sg13g2_xnor2_1
X_4668_ _1482_ _1479_ _1481_ VPWR VGND sg13g2_nand2_1
X_3619_ VGND VPWR _0478_ _0476_ _0436_ sg13g2_or2_1
X_6407_ net1073 VGND VPWR net214 mac2.sum_lvl1_ff\[40\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_4599_ _1415_ _1414_ _1413_ VPWR VGND sg13g2_nand2b_1
X_6338_ net1020 VGND VPWR net411 mac1.total_sum\[15\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_6269_ net1026 VGND VPWR net211 mac2.sum_lvl1_ff\[82\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_44_32 VPWR VGND sg13g2_fill_2
XFILLER_25_550 VPWR VGND sg13g2_fill_2
XFILLER_8_226 VPWR VGND sg13g2_fill_2
XFILLER_8_248 VPWR VGND sg13g2_fill_1
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_48_653 VPWR VGND sg13g2_fill_1
XFILLER_35_314 VPWR VGND sg13g2_fill_1
XFILLER_35_325 VPWR VGND sg13g2_fill_2
X_3970_ _0765_ _0812_ _0814_ VPWR VGND sg13g2_and2_1
X_5640_ _2351_ _2352_ net22 VPWR VGND sg13g2_nor2b_1
XFILLER_31_575 VPWR VGND sg13g2_decap_4
X_5571_ _2299_ mac2.sum_lvl3_ff\[34\] net347 VPWR VGND sg13g2_nand2_1
X_4522_ _1344_ _1327_ _1343_ VPWR VGND sg13g2_xnor2_1
Xhold226 _0000_ VPWR VGND net266 sg13g2_dlygate4sd3_1
Xhold215 mac2.products_ff\[140\] VPWR VGND net255 sg13g2_dlygate4sd3_1
Xhold204 mac2.sum_lvl1_ff\[1\] VPWR VGND net244 sg13g2_dlygate4sd3_1
X_4453_ _1278_ net859 net803 VPWR VGND sg13g2_nand2_1
Xhold248 DP_4.matrix\[73\] VPWR VGND net288 sg13g2_dlygate4sd3_1
X_3404_ _0269_ net992 net928 VPWR VGND sg13g2_nand2_1
Xhold237 DP_2.matrix\[72\] VPWR VGND net277 sg13g2_dlygate4sd3_1
Xhold259 DP_1.matrix\[72\] VPWR VGND net299 sg13g2_dlygate4sd3_1
X_4384_ VGND VPWR _1211_ _1209_ _1170_ sg13g2_or2_1
X_6123_ net1077 VGND VPWR _0235_ DP_3.matrix\[43\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3335_ _2922_ _2885_ _2920_ VPWR VGND sg13g2_xnor2_1
X_3266_ _2838_ _2831_ _2799_ _2855_ VPWR VGND sg13g2_a21o_1
X_6054_ net1039 VGND VPWR _0189_ DP_1.matrix\[73\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_5005_ _1801_ _1802_ _1796_ _1804_ VPWR VGND sg13g2_nand3_1
XFILLER_39_642 VPWR VGND sg13g2_fill_2
X_3197_ _2787_ _2779_ _2788_ VPWR VGND sg13g2_nor2b_1
X_5907_ _2581_ VPWR _0249_ VGND net761 _2582_ sg13g2_o21ai_1
X_5838_ net983 net756 _2538_ VPWR VGND sg13g2_nor2_1
X_5769_ _2473_ VPWR _2476_ VGND _2474_ _2475_ sg13g2_o21ai_1
XFILLER_2_936 VPWR VGND sg13g2_decap_8
XFILLER_45_601 VPWR VGND sg13g2_fill_1
X_3120_ _2709_ _2710_ _2712_ _2713_ VPWR VGND sg13g2_or3_1
XFILLER_49_940 VPWR VGND sg13g2_decap_8
X_3051_ _2646_ net946 net904 net949 net898 VPWR VGND sg13g2_a22oi_1
XFILLER_35_133 VPWR VGND sg13g2_fill_1
X_3953_ _0760_ VPWR _0797_ VGND _0718_ _0761_ sg13g2_o21ai_1
XFILLER_16_391 VPWR VGND sg13g2_fill_1
X_3884_ DP_2.matrix\[36\] net919 net963 net962 _0730_ VPWR VGND sg13g2_and4_1
X_5623_ _2338_ _2336_ net19 VPWR VGND sg13g2_xor2_1
XFILLER_8_590 VPWR VGND sg13g2_decap_4
X_5554_ VGND VPWR _2285_ mac2.sum_lvl3_ff\[11\] net423 sg13g2_or2_1
X_4505_ _1328_ net803 net1000 VPWR VGND sg13g2_nand2_1
X_5485_ VGND VPWR _2226_ _2228_ _2232_ _2225_ sg13g2_a21oi_1
X_4436_ _1262_ _1241_ _1261_ VPWR VGND sg13g2_xnor2_1
X_4367_ _1195_ _1165_ _1194_ VPWR VGND sg13g2_nand2_1
X_6106_ net1066 VGND VPWR net68 mac1.sum_lvl1_ff\[3\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3318_ _2904_ _2903_ _2906_ VPWR VGND sg13g2_xor2_1
X_4298_ _1127_ _1120_ _1126_ VPWR VGND sg13g2_nand2_1
X_3249_ _2839_ _2831_ _2838_ VPWR VGND sg13g2_xnor2_1
X_6037_ net1044 VGND VPWR _0174_ DP_1.matrix\[2\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_26_122 VPWR VGND sg13g2_fill_2
XFILLER_26_133 VPWR VGND sg13g2_fill_2
XFILLER_25_67 VPWR VGND sg13g2_fill_1
XFILLER_6_505 VPWR VGND sg13g2_fill_2
XFILLER_9_2 VPWR VGND sg13g2_fill_1
XFILLER_1_243 VPWR VGND sg13g2_fill_1
XFILLER_49_225 VPWR VGND sg13g2_fill_1
XFILLER_2_27 VPWR VGND sg13g2_fill_2
XFILLER_46_910 VPWR VGND sg13g2_decap_8
XFILLER_46_987 VPWR VGND sg13g2_decap_8
XFILLER_40_180 VPWR VGND sg13g2_fill_2
X_5270_ _2061_ net841 net994 VPWR VGND sg13g2_nand2_1
X_4221_ _1052_ _1050_ _1051_ VPWR VGND sg13g2_nand2b_1
X_4152_ _0986_ _0983_ _0987_ VPWR VGND sg13g2_xor2_1
X_3103_ _2696_ net887 net958 net889 net957 VPWR VGND sg13g2_a22oi_1
X_4083_ VGND VPWR _0874_ _0893_ _0924_ _0895_ sg13g2_a21oi_1
XFILLER_28_409 VPWR VGND sg13g2_fill_1
XFILLER_49_792 VPWR VGND sg13g2_decap_4
X_3034_ _2629_ _2619_ _2630_ VPWR VGND sg13g2_xor2_1
XFILLER_37_965 VPWR VGND sg13g2_decap_8
XFILLER_36_486 VPWR VGND sg13g2_fill_2
XFILLER_24_648 VPWR VGND sg13g2_decap_8
X_4985_ _1784_ _1776_ _1780_ VPWR VGND sg13g2_nand2_1
X_3936_ _0770_ _0778_ _0780_ _0781_ VPWR VGND sg13g2_or3_1
XFILLER_32_670 VPWR VGND sg13g2_fill_1
X_3867_ _0713_ _0712_ _0123_ VPWR VGND sg13g2_xor2_1
X_3798_ _0645_ _0646_ _0640_ _0647_ VPWR VGND sg13g2_nand3_1
X_5606_ _2325_ mac1.total_sum\[7\] mac2.total_sum\[7\] VPWR VGND sg13g2_nand2_1
X_5537_ _2271_ VPWR _2272_ VGND _2265_ _2268_ sg13g2_o21ai_1
XFILLER_11_69 VPWR VGND sg13g2_fill_2
X_5468_ _2217_ _2218_ _0045_ VPWR VGND sg13g2_and2_1
X_4419_ VGND VPWR _1245_ _1244_ _1220_ sg13g2_or2_1
X_5399_ VGND VPWR _2160_ _2162_ _2165_ net406 sg13g2_a21oi_1
XFILLER_28_965 VPWR VGND sg13g2_decap_8
XFILLER_43_913 VPWR VGND sg13g2_decap_8
XFILLER_14_103 VPWR VGND sg13g2_fill_1
Xheichips25_SDR_33 VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_7_836 VPWR VGND sg13g2_fill_1
XFILLER_2_596 VPWR VGND sg13g2_fill_2
XFILLER_19_987 VPWR VGND sg13g2_decap_8
XFILLER_33_401 VPWR VGND sg13g2_fill_2
XFILLER_45_283 VPWR VGND sg13g2_fill_2
XFILLER_34_968 VPWR VGND sg13g2_decap_8
X_4770_ _1581_ _1574_ _1580_ VPWR VGND sg13g2_xnor2_1
X_3721_ _0538_ _0576_ _0577_ VPWR VGND sg13g2_nor2_1
X_3652_ _0510_ DP_2.matrix\[3\] net1011 VPWR VGND sg13g2_nand2_1
X_6440_ net1057 VGND VPWR net139 mac2.sum_lvl2_ff\[19\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3583_ _0412_ VPWR _0443_ VGND _0403_ _0413_ sg13g2_o21ai_1
X_6371_ net1050 VGND VPWR _0089_ mac2.products_ff\[136\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5322_ _2105_ net499 mac1.sum_lvl2_ff\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_47_0 VPWR VGND sg13g2_decap_4
X_5253_ _2045_ _2009_ _2043_ VPWR VGND sg13g2_xnor2_1
X_5184_ _1961_ _1955_ _1923_ _1978_ VPWR VGND sg13g2_a21o_1
X_4204_ _1036_ _1029_ _1034_ _1035_ VPWR VGND sg13g2_and3_1
X_4135_ VGND VPWR _0956_ _0972_ _0973_ _0971_ sg13g2_a21oi_1
X_4066_ _0878_ VPWR _0907_ VGND _0876_ _0879_ sg13g2_o21ai_1
XFILLER_37_751 VPWR VGND sg13g2_fill_2
X_3017_ _2614_ _2602_ _2612_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_927 VPWR VGND sg13g2_decap_8
X_4968_ _1768_ net845 net798 net847 net795 VPWR VGND sg13g2_a22oi_1
X_4899_ _1692_ _1705_ _1706_ VPWR VGND sg13g2_nor2_1
X_3919_ _0764_ net971 net910 VPWR VGND sg13g2_nand2_1
XFILLER_47_76 VPWR VGND sg13g2_fill_1
XFILLER_16_913 VPWR VGND sg13g2_decap_8
XFILLER_43_787 VPWR VGND sg13g2_decap_8
XFILLER_31_927 VPWR VGND sg13g2_decap_8
XFILLER_10_150 VPWR VGND sg13g2_fill_2
XFILLER_10_172 VPWR VGND sg13g2_fill_1
X_5940_ net916 _0206_ VPWR VGND sg13g2_buf_1
XFILLER_33_220 VPWR VGND sg13g2_fill_1
X_5871_ _2467_ _2462_ _2559_ VPWR VGND sg13g2_xor2_1
X_4822_ _1599_ _1630_ _1597_ _1632_ VPWR VGND sg13g2_nand3_1
X_4753_ _1563_ _1531_ _1565_ VPWR VGND sg13g2_xor2_1
X_3704_ VGND VPWR _0500_ _0533_ _0561_ _0532_ sg13g2_a21oi_1
X_6423_ net1027 VGND VPWR net4 DP_1.I_range.out_data\[6\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_4684_ _1470_ VPWR _1497_ VGND _1461_ _1471_ sg13g2_o21ai_1
X_3635_ _0492_ _0484_ _0494_ VPWR VGND sg13g2_xor2_1
X_6354_ net1092 VGND VPWR _0144_ mac2.products_ff\[15\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3566_ _0424_ _0423_ _0425_ _0427_ VPWR VGND sg13g2_a21o_1
X_5305_ _2092_ mac1.sum_lvl2_ff\[22\] mac1.sum_lvl2_ff\[3\] VPWR VGND sg13g2_nand2_1
X_3497_ _0359_ _0321_ _0357_ VPWR VGND sg13g2_xnor2_1
X_6285_ net1020 VGND VPWR net123 mac1.sum_lvl3_ff\[30\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_5236_ _2027_ _2028_ _2029_ VPWR VGND sg13g2_nor2_1
XFILLER_25_1022 VPWR VGND sg13g2_decap_8
X_5167_ _1962_ _1955_ _1961_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_526 VPWR VGND sg13g2_fill_2
X_4118_ _0946_ _0948_ _0957_ VPWR VGND sg13g2_and2_1
X_5098_ _1848_ VPWR _1895_ VGND _1787_ _1849_ sg13g2_o21ai_1
X_4049_ _0889_ _0882_ _0891_ VPWR VGND sg13g2_xor2_1
XFILLER_37_570 VPWR VGND sg13g2_decap_4
XFILLER_24_264 VPWR VGND sg13g2_fill_1
XFILLER_32_1004 VPWR VGND sg13g2_decap_8
XFILLER_40_757 VPWR VGND sg13g2_fill_1
Xhold8 mac2.sum_lvl2_ff\[51\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_35_529 VPWR VGND sg13g2_fill_2
XFILLER_8_931 VPWR VGND sg13g2_decap_8
XFILLER_12_971 VPWR VGND sg13g2_decap_8
XFILLER_7_463 VPWR VGND sg13g2_fill_1
Xhold408 mac2.sum_lvl2_ff\[5\] VPWR VGND net448 sg13g2_dlygate4sd3_1
X_3420_ _0283_ _0282_ _0285_ VPWR VGND sg13g2_xor2_1
Xhold419 _2269_ VPWR VGND net459 sg13g2_dlygate4sd3_1
X_3351_ _2926_ _2928_ _2937_ VPWR VGND sg13g2_and2_1
X_6070_ net1015 VGND VPWR _0102_ mac1.products_ff\[143\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3282_ _2870_ _2862_ _2871_ VPWR VGND sg13g2_nor2b_1
X_5021_ _1819_ net852 net781 VPWR VGND sg13g2_nand2_1
XFILLER_38_356 VPWR VGND sg13g2_fill_2
XFILLER_47_890 VPWR VGND sg13g2_decap_8
X_5923_ net976 _0181_ VPWR VGND sg13g2_buf_1
X_5854_ VGND VPWR net757 _2548_ _0198_ _2546_ sg13g2_a21oi_1
XFILLER_34_584 VPWR VGND sg13g2_fill_2
X_4805_ _1615_ _1609_ _1614_ VPWR VGND sg13g2_xnor2_1
X_5785_ VGND VPWR _2489_ _2490_ _0166_ _2491_ sg13g2_a21oi_1
X_2997_ _2594_ _2595_ _0065_ VPWR VGND sg13g2_nor2_1
X_4736_ _1499_ _1546_ _1548_ VPWR VGND sg13g2_and2_1
X_4667_ _1478_ _1477_ _1448_ _1481_ VPWR VGND sg13g2_a21o_1
X_3618_ _0477_ net986 net926 VPWR VGND sg13g2_nand2_1
X_6406_ net1072 VGND VPWR net79 mac2.sum_lvl1_ff\[39\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_6337_ net1018 VGND VPWR net375 mac1.total_sum\[14\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_4598_ _1386_ VPWR _1414_ VGND _1410_ _1411_ sg13g2_o21ai_1
X_3549_ _0405_ VPWR _0410_ VGND _0406_ _0408_ sg13g2_o21ai_1
X_6268_ net1028 VGND VPWR net54 mac2.sum_lvl1_ff\[81\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_5219_ _1981_ VPWR _2012_ VGND _1979_ _1982_ sg13g2_o21ai_1
X_6199_ net1068 VGND VPWR net160 mac1.sum_lvl2_ff\[23\] clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_12_234 VPWR VGND sg13g2_fill_2
XFILLER_12_256 VPWR VGND sg13g2_fill_2
XFILLER_12_289 VPWR VGND sg13g2_fill_2
XFILLER_4_433 VPWR VGND sg13g2_fill_1
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_499 VPWR VGND sg13g2_fill_1
XFILLER_0_672 VPWR VGND sg13g2_fill_2
XFILLER_47_142 VPWR VGND sg13g2_fill_2
XFILLER_44_893 VPWR VGND sg13g2_decap_8
XFILLER_31_598 VPWR VGND sg13g2_fill_1
X_5570_ VGND VPWR mac2.sum_lvl3_ff\[33\] mac2.sum_lvl3_ff\[13\] _2298_ _2296_ sg13g2_a21oi_1
X_4521_ _1343_ net856 DP_4.matrix\[44\] VPWR VGND sg13g2_nand2_1
Xhold216 mac2.sum_lvl2_ff\[38\] VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold205 mac2.products_ff\[142\] VPWR VGND net245 sg13g2_dlygate4sd3_1
X_4452_ _1277_ net858 net801 VPWR VGND sg13g2_nand2_1
X_3403_ _0268_ net928 net993 net929 net992 VPWR VGND sg13g2_a22oi_1
Xhold238 DP_1.matrix\[78\] VPWR VGND net278 sg13g2_dlygate4sd3_1
Xhold227 mac2.sum_lvl2_ff\[0\] VPWR VGND net267 sg13g2_dlygate4sd3_1
Xhold249 _1717_ VPWR VGND net289 sg13g2_dlygate4sd3_1
X_4383_ _1210_ net864 net804 VPWR VGND sg13g2_nand2_1
X_6122_ net1092 VGND VPWR _0234_ DP_3.matrix\[42\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3334_ _2885_ _2920_ _2921_ VPWR VGND sg13g2_nor2b_1
X_6053_ net1040 VGND VPWR _0188_ DP_1.matrix\[72\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_3265_ _2840_ VPWR _2854_ VGND _2829_ _2841_ sg13g2_o21ai_1
XFILLER_22_1025 VPWR VGND sg13g2_decap_4
X_5004_ _1803_ _1796_ _1801_ _1802_ VPWR VGND sg13g2_and3_1
X_3196_ _2787_ _2780_ _2786_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_698 VPWR VGND sg13g2_fill_2
X_5906_ _2515_ _2497_ _2582_ VPWR VGND sg13g2_xor2_1
X_5837_ VGND VPWR net753 _2537_ _0176_ _2536_ sg13g2_a21oi_1
X_5768_ net767 VPWR _2475_ VGND net878 net778 sg13g2_o21ai_1
X_4719_ _1494_ VPWR _1531_ VGND _1452_ _1495_ sg13g2_o21ai_1
X_5699_ _2375_ _2407_ _2408_ VPWR VGND sg13g2_nor2_1
XFILLER_2_915 VPWR VGND sg13g2_decap_8
XFILLER_1_403 VPWR VGND sg13g2_fill_2
XFILLER_44_112 VPWR VGND sg13g2_fill_1
XFILLER_17_337 VPWR VGND sg13g2_fill_1
XFILLER_41_885 VPWR VGND sg13g2_decap_8
XFILLER_45_1014 VPWR VGND sg13g2_decap_8
X_3050_ net901 net949 net904 _2645_ VPWR VGND net946 sg13g2_nand4_1
XFILLER_49_996 VPWR VGND sg13g2_decap_8
XFILLER_35_123 VPWR VGND sg13g2_fill_1
XFILLER_17_882 VPWR VGND sg13g2_fill_2
X_3952_ _0125_ _0751_ _0795_ VPWR VGND sg13g2_xnor2_1
X_3883_ _0729_ net916 net966 VPWR VGND sg13g2_nand2_1
XFILLER_32_885 VPWR VGND sg13g2_decap_8
X_5622_ _2333_ _2337_ _2338_ VPWR VGND sg13g2_nor2_1
X_5553_ net423 mac2.sum_lvl3_ff\[11\] _2284_ VPWR VGND sg13g2_and2_1
X_4504_ _1327_ net801 net1000 VPWR VGND sg13g2_nand2_1
X_5484_ _2229_ _2230_ _2231_ VPWR VGND sg13g2_nor2b_1
X_4435_ _1259_ _1248_ _1261_ VPWR VGND sg13g2_xor2_1
X_4366_ _1193_ _1176_ _1194_ VPWR VGND sg13g2_xor2_1
X_3317_ VGND VPWR _2905_ _2904_ _2903_ sg13g2_or2_1
X_6105_ net1060 VGND VPWR _0223_ DP_3.matrix\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4297_ _1126_ _1121_ _1124_ VPWR VGND sg13g2_xnor2_1
X_3248_ _2836_ _2837_ _2838_ VPWR VGND sg13g2_nor2b_1
X_6036_ net1044 VGND VPWR _0173_ DP_1.matrix\[1\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3179_ _2768_ _2769_ _2700_ _2771_ VPWR VGND sg13g2_nand3_1
XFILLER_26_112 VPWR VGND sg13g2_fill_1
XFILLER_39_473 VPWR VGND sg13g2_fill_2
XFILLER_41_12 VPWR VGND sg13g2_fill_1
XFILLER_45_410 VPWR VGND sg13g2_fill_1
XFILLER_17_101 VPWR VGND sg13g2_fill_1
XFILLER_46_966 VPWR VGND sg13g2_decap_8
XFILLER_17_167 VPWR VGND sg13g2_fill_2
XFILLER_12_1013 VPWR VGND sg13g2_decap_8
XFILLER_5_561 VPWR VGND sg13g2_fill_1
X_4220_ _1051_ net871 net803 VPWR VGND sg13g2_nand2_1
X_4151_ _0984_ _0985_ _0986_ VPWR VGND sg13g2_nor2_1
X_3102_ _2672_ VPWR _2695_ VGND _2637_ _2670_ sg13g2_o21ai_1
X_4082_ _0923_ _0901_ _0922_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_771 VPWR VGND sg13g2_decap_8
X_3033_ _2629_ _2627_ _2628_ VPWR VGND sg13g2_nand2_1
XFILLER_37_944 VPWR VGND sg13g2_decap_8
X_4984_ _0149_ _1756_ _1783_ VPWR VGND sg13g2_xnor2_1
X_3935_ VGND VPWR _0776_ _0777_ _0780_ _0771_ sg13g2_a21oi_1
XFILLER_32_693 VPWR VGND sg13g2_decap_4
X_3866_ VGND VPWR _0654_ _0680_ _0713_ _0679_ sg13g2_a21oi_1
X_5605_ _2323_ _2324_ net31 VPWR VGND sg13g2_nor2b_1
X_3797_ _0641_ VPWR _0646_ VGND _0642_ _0644_ sg13g2_o21ai_1
X_5536_ net539 net436 _2271_ VPWR VGND sg13g2_xor2_1
X_5467_ _2210_ _2213_ _2216_ _2218_ VPWR VGND sg13g2_or3_1
X_4418_ _1244_ net810 net1000 VPWR VGND sg13g2_nand2_1
X_5398_ _2164_ mac1.sum_lvl3_ff\[28\] net405 VPWR VGND sg13g2_xnor2_1
X_4349_ _1146_ VPWR _1177_ VGND _1137_ _1147_ sg13g2_o21ai_1
X_6019_ net1083 VGND VPWR _0119_ mac1.products_ff\[80\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_27_410 VPWR VGND sg13g2_fill_2
XFILLER_28_944 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_43_969 VPWR VGND sg13g2_decap_8
XFILLER_35_1013 VPWR VGND sg13g2_decap_8
Xheichips25_SDR_34 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_11_877 VPWR VGND sg13g2_fill_1
Xfanout890 net891 net890 VPWR VGND sg13g2_buf_8
XFILLER_19_966 VPWR VGND sg13g2_decap_8
XFILLER_33_424 VPWR VGND sg13g2_fill_1
XFILLER_34_947 VPWR VGND sg13g2_decap_8
XFILLER_33_468 VPWR VGND sg13g2_fill_1
XFILLER_42_980 VPWR VGND sg13g2_decap_8
X_3720_ _0576_ _0567_ _0575_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_130 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_40_clk clknet_4_12_0_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ _0509_ DP_2.matrix\[5\] net982 VPWR VGND sg13g2_nand2_1
X_6370_ net1093 VGND VPWR _0133_ mac2.products_ff\[83\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3582_ _0440_ _0432_ _0442_ VPWR VGND sg13g2_xor2_1
X_5321_ _2103_ net516 _0012_ VPWR VGND sg13g2_nor2b_2
X_5252_ _2009_ _2043_ _2044_ VPWR VGND sg13g2_nor2b_1
X_4203_ _1030_ VPWR _1035_ VGND _1031_ _1033_ sg13g2_o21ai_1
X_5183_ _1963_ VPWR _1977_ VGND _1953_ _1964_ sg13g2_o21ai_1
X_4134_ _0972_ _0956_ _0121_ VPWR VGND sg13g2_xor2_1
X_4065_ _0886_ VPWR _0906_ VGND _0884_ _0887_ sg13g2_o21ai_1
X_3016_ _2613_ _2612_ _2602_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_903 VPWR VGND sg13g2_decap_4
XFILLER_19_1008 VPWR VGND sg13g2_decap_8
XFILLER_40_906 VPWR VGND sg13g2_decap_8
X_4967_ net795 net846 net798 _1767_ VPWR VGND net844 sg13g2_nand4_1
X_4898_ _1703_ _1693_ _1705_ VPWR VGND sg13g2_xor2_1
X_3918_ _0736_ VPWR _0763_ VGND _0727_ _0737_ sg13g2_o21ai_1
Xclkbuf_leaf_31_clk clknet_4_13_0_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_3849_ net922 net921 net967 net965 _0696_ VPWR VGND sg13g2_and4_1
X_5519_ _2258_ mac2.sum_lvl3_ff\[23\] net487 VPWR VGND sg13g2_xnor2_1
XFILLER_43_744 VPWR VGND sg13g2_fill_2
XFILLER_43_722 VPWR VGND sg13g2_fill_1
XFILLER_43_755 VPWR VGND sg13g2_fill_2
XFILLER_31_906 VPWR VGND sg13g2_decap_8
XFILLER_8_27 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_22_clk clknet_4_5_0_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_6_177 VPWR VGND sg13g2_fill_1
XFILLER_3_862 VPWR VGND sg13g2_fill_2
XFILLER_2_350 VPWR VGND sg13g2_fill_1
X_5870_ _0220_ net886 net758 VPWR VGND sg13g2_xnor2_1
XFILLER_22_917 VPWR VGND sg13g2_fill_1
X_4821_ VGND VPWR _1597_ _1599_ _1631_ _1630_ sg13g2_a21oi_1
XFILLER_15_980 VPWR VGND sg13g2_decap_8
XFILLER_21_438 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_13_clk clknet_4_6_0_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4752_ _1564_ _1531_ _1563_ VPWR VGND sg13g2_nand2b_1
X_3703_ _0558_ _0557_ _0560_ VPWR VGND sg13g2_xor2_1
XFILLER_30_983 VPWR VGND sg13g2_decap_8
X_4683_ _1496_ _1452_ _1495_ VPWR VGND sg13g2_xnor2_1
X_3634_ _0493_ _0484_ _0492_ VPWR VGND sg13g2_nand2b_1
X_6422_ net1027 VGND VPWR DP_1.I_range.data_plus_4\[6\] DP_1.I_range.out_data\[5\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_6353_ net1092 VGND VPWR _0143_ mac2.products_ff\[14\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3565_ _0424_ _0425_ _0423_ _0426_ VPWR VGND sg13g2_nand3_1
X_5304_ VGND VPWR _2088_ _2090_ _2091_ _2089_ sg13g2_a21oi_1
X_3496_ VGND VPWR _0358_ _0356_ _0322_ sg13g2_or2_1
X_6284_ net1020 VGND VPWR net58 mac1.sum_lvl3_ff\[29\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_5235_ VGND VPWR _1977_ _1998_ _2028_ _2000_ sg13g2_a21oi_1
XFILLER_25_1001 VPWR VGND sg13g2_decap_8
X_5166_ _1960_ _1956_ _1961_ VPWR VGND sg13g2_xor2_1
X_4117_ _0954_ _0930_ _0955_ _0956_ VPWR VGND sg13g2_a21o_1
X_5097_ _1891_ _1892_ _1822_ _1894_ VPWR VGND sg13g2_nand3_1
X_4048_ _0889_ _0882_ _0890_ VPWR VGND sg13g2_nor2b_1
X_5999_ net1070 VGND VPWR _0114_ mac1.products_ff\[8\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_21_983 VPWR VGND sg13g2_decap_8
XFILLER_33_79 VPWR VGND sg13g2_fill_1
XFILLER_4_659 VPWR VGND sg13g2_fill_2
XFILLER_3_125 VPWR VGND sg13g2_fill_1
XFILLER_47_313 VPWR VGND sg13g2_fill_1
Xhold9 mac1.sum_lvl1_ff\[11\] VPWR VGND net49 sg13g2_dlygate4sd3_1
XFILLER_47_357 VPWR VGND sg13g2_fill_1
XFILLER_12_950 VPWR VGND sg13g2_decap_8
XFILLER_8_987 VPWR VGND sg13g2_decap_8
Xhold409 _2209_ VPWR VGND net449 sg13g2_dlygate4sd3_1
X_3350_ _2934_ _2910_ _2935_ _2936_ VPWR VGND sg13g2_a21o_1
X_3281_ _2870_ _2863_ _2869_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_4 VPWR VGND sg13g2_fill_1
X_5020_ _1818_ net781 net854 net783 net852 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_38_335 VPWR VGND sg13g2_fill_2
XFILLER_0_1025 VPWR VGND sg13g2_decap_4
X_5922_ net281 _0180_ VPWR VGND sg13g2_buf_1
X_5853_ _2548_ _2429_ _2547_ VPWR VGND sg13g2_nand2_1
X_5784_ _2451_ _2490_ _2491_ VPWR VGND sg13g2_nor2_1
X_4804_ _1613_ _1610_ _1614_ VPWR VGND sg13g2_xor2_1
X_4735_ VGND VPWR _1547_ _1546_ _1499_ sg13g2_or2_1
X_2996_ _2595_ net898 net958 net956 net903 VPWR VGND sg13g2_a22oi_1
X_4666_ VGND VPWR _1477_ _1478_ _1480_ _1448_ sg13g2_a21oi_1
X_3617_ _0476_ net986 net925 VPWR VGND sg13g2_nand2_1
X_6405_ net1059 VGND VPWR net203 mac2.sum_lvl1_ff\[38\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4597_ _1386_ _1410_ _1411_ _1413_ VPWR VGND sg13g2_nor3_1
X_3548_ _0405_ _0406_ _0408_ _0409_ VPWR VGND sg13g2_or3_1
X_6336_ net1017 VGND VPWR net343 mac1.total_sum\[13\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3479_ _0342_ _0318_ _0341_ VPWR VGND sg13g2_xnor2_1
X_6267_ net1028 VGND VPWR net132 mac2.sum_lvl1_ff\[80\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_6198_ net1067 VGND VPWR net116 mac1.sum_lvl2_ff\[22\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_5218_ _1992_ VPWR _2011_ VGND _1946_ _1990_ sg13g2_o21ai_1
XFILLER_28_46 VPWR VGND sg13g2_fill_2
XFILLER_29_324 VPWR VGND sg13g2_fill_2
X_5149_ _1917_ VPWR _1944_ VGND _1914_ _1918_ sg13g2_o21ai_1
XFILLER_37_390 VPWR VGND sg13g2_fill_2
XFILLER_40_511 VPWR VGND sg13g2_fill_1
XFILLER_13_769 VPWR VGND sg13g2_fill_1
XFILLER_40_533 VPWR VGND sg13g2_fill_2
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_35_327 VPWR VGND sg13g2_fill_1
XFILLER_16_552 VPWR VGND sg13g2_decap_4
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
X_4520_ _1330_ VPWR _1342_ VGND _1304_ _1327_ sg13g2_o21ai_1
XFILLER_8_773 VPWR VGND sg13g2_fill_2
X_4451_ _1276_ net864 net995 VPWR VGND sg13g2_nand2_1
XFILLER_7_261 VPWR VGND sg13g2_fill_2
Xhold217 mac1.products_ff\[79\] VPWR VGND net257 sg13g2_dlygate4sd3_1
Xhold206 mac2.sum_lvl1_ff\[42\] VPWR VGND net246 sg13g2_dlygate4sd3_1
X_3402_ _0072_ _2968_ _2981_ VPWR VGND sg13g2_xnor2_1
Xhold228 _0032_ VPWR VGND net268 sg13g2_dlygate4sd3_1
Xhold239 DP_3.matrix\[72\] VPWR VGND net279 sg13g2_dlygate4sd3_1
X_4382_ _1209_ net864 net802 VPWR VGND sg13g2_nand2_1
X_6121_ net1070 VGND VPWR net61 mac1.sum_lvl1_ff\[8\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_3333_ _2920_ _2915_ _2918_ VPWR VGND sg13g2_xnor2_1
X_6052_ net1039 VGND VPWR _0065_ mac1.products_ff\[137\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_3264_ _2826_ _2820_ _2828_ _2853_ VPWR VGND sg13g2_a21o_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
XFILLER_22_1004 VPWR VGND sg13g2_decap_8
X_5003_ _1797_ VPWR _1802_ VGND _1798_ _1800_ sg13g2_o21ai_1
X_3195_ _2785_ _2781_ _2786_ VPWR VGND sg13g2_xor2_1
X_5905_ _2581_ net822 net761 VPWR VGND sg13g2_nand2_1
XFILLER_35_894 VPWR VGND sg13g2_decap_8
X_5836_ _2399_ _2395_ _2537_ VPWR VGND sg13g2_xor2_1
X_5767_ net863 net779 _2474_ VPWR VGND sg13g2_nor2_1
X_5698_ net755 VPWR _2407_ VGND _2404_ _2406_ sg13g2_o21ai_1
X_4718_ _0147_ _1485_ _1529_ VPWR VGND sg13g2_xnor2_1
X_4649_ _1463_ net827 net877 VPWR VGND sg13g2_nand2_1
X_6319_ net1029 VGND VPWR net82 mac2.sum_lvl3_ff\[32\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_45_636 VPWR VGND sg13g2_fill_1
XFILLER_25_371 VPWR VGND sg13g2_fill_1
XFILLER_26_894 VPWR VGND sg13g2_decap_8
XFILLER_13_555 VPWR VGND sg13g2_fill_1
XFILLER_41_864 VPWR VGND sg13g2_decap_8
XFILLER_49_975 VPWR VGND sg13g2_decap_8
XFILLER_48_474 VPWR VGND sg13g2_fill_2
XFILLER_35_146 VPWR VGND sg13g2_fill_1
X_3951_ _0750_ _0795_ _0749_ _0796_ VPWR VGND sg13g2_nand3_1
XFILLER_44_691 VPWR VGND sg13g2_fill_1
X_3882_ _0697_ VPWR _0728_ VGND _0695_ _0698_ sg13g2_o21ai_1
X_5621_ VPWR VGND mac2.total_sum\[9\] _2330_ mac1.total_sum\[9\] mac1.total_sum\[8\]
+ _2337_ mac2.total_sum\[8\] sg13g2_a221oi_1
X_5552_ _2283_ net381 _0049_ VPWR VGND sg13g2_xor2_1
X_4503_ _1326_ net858 net995 VPWR VGND sg13g2_nand2_1
X_5483_ VGND VPWR _2230_ mac2.sum_lvl2_ff\[11\] mac2.sum_lvl2_ff\[30\] sg13g2_or2_1
X_4434_ _1248_ _1259_ _1260_ VPWR VGND sg13g2_nor2_1
X_4365_ _1193_ _1177_ _1191_ VPWR VGND sg13g2_xnor2_1
X_3316_ VGND VPWR _2854_ _2874_ _2904_ _2876_ sg13g2_a21oi_1
X_6104_ net1060 VGND VPWR _0222_ DP_3.matrix\[2\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6035_ net1044 VGND VPWR _0172_ DP_1.matrix\[0\] clknet_leaf_56_clk sg13g2_dfrbpq_2
X_4296_ _1125_ _1124_ _1121_ VPWR VGND sg13g2_nand2b_1
X_3247_ _2832_ VPWR _2837_ VGND _2834_ _2835_ sg13g2_o21ai_1
X_3178_ _2769_ _2768_ _2700_ _2770_ VPWR VGND sg13g2_a21o_1
XFILLER_27_669 VPWR VGND sg13g2_fill_1
XFILLER_22_341 VPWR VGND sg13g2_fill_1
X_5819_ net760 _2493_ _2525_ VPWR VGND sg13g2_nor2_1
XFILLER_46_945 VPWR VGND sg13g2_decap_8
XFILLER_18_625 VPWR VGND sg13g2_decap_4
XFILLER_33_606 VPWR VGND sg13g2_fill_1
XFILLER_33_628 VPWR VGND sg13g2_fill_1
XFILLER_13_385 VPWR VGND sg13g2_fill_2
X_4150_ _0985_ net867 net819 net440 net869 VPWR VGND sg13g2_a22oi_1
X_3101_ _2686_ VPWR _2694_ VGND _2666_ _2687_ sg13g2_o21ai_1
XFILLER_49_750 VPWR VGND sg13g2_decap_8
X_4081_ _0922_ _0919_ _0920_ VPWR VGND sg13g2_xnor2_1
X_3032_ _2626_ _2625_ _2620_ _2628_ VPWR VGND sg13g2_a21o_1
XFILLER_37_923 VPWR VGND sg13g2_decap_8
X_4983_ _1783_ _1782_ _1781_ VPWR VGND sg13g2_nand2b_1
X_3934_ _0776_ _0777_ _0771_ _0779_ VPWR VGND sg13g2_nand3_1
X_3865_ _0710_ _0682_ _0712_ VPWR VGND sg13g2_xor2_1
XFILLER_20_812 VPWR VGND sg13g2_fill_1
X_5604_ _2321_ VPWR _2324_ VGND _2318_ _2322_ sg13g2_o21ai_1
XFILLER_20_856 VPWR VGND sg13g2_fill_2
X_3796_ _0641_ _0642_ _0644_ _0645_ VPWR VGND sg13g2_or3_1
X_5535_ _2270_ net436 mac2.sum_lvl3_ff\[7\] VPWR VGND sg13g2_nand2_1
X_5466_ _2216_ VPWR _2217_ VGND _2210_ _2213_ sg13g2_o21ai_1
X_4417_ _1243_ net805 net859 VPWR VGND sg13g2_nand2_1
X_5397_ net520 _2163_ _0029_ VPWR VGND sg13g2_and2_1
XFILLER_28_1021 VPWR VGND sg13g2_decap_8
X_4348_ _1174_ _1166_ _1176_ VPWR VGND sg13g2_xor2_1
X_4279_ VGND VPWR _1105_ _1106_ _1109_ _1089_ sg13g2_a21oi_1
X_6018_ net1086 VGND VPWR _0118_ mac1.products_ff\[79\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_28_923 VPWR VGND sg13g2_decap_8
XFILLER_27_466 VPWR VGND sg13g2_decap_8
XFILLER_36_79 VPWR VGND sg13g2_fill_2
XFILLER_43_948 VPWR VGND sg13g2_decap_8
XFILLER_42_469 VPWR VGND sg13g2_decap_4
XFILLER_11_812 VPWR VGND sg13g2_fill_1
XFILLER_23_683 VPWR VGND sg13g2_fill_2
Xheichips25_SDR_35 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_2_598 VPWR VGND sg13g2_fill_1
XFILLER_38_709 VPWR VGND sg13g2_fill_2
Xfanout891 net357 net891 VPWR VGND sg13g2_buf_1
XFILLER_19_923 VPWR VGND sg13g2_decap_8
Xfanout880 net881 net880 VPWR VGND sg13g2_buf_8
XFILLER_34_926 VPWR VGND sg13g2_decap_8
XFILLER_9_153 VPWR VGND sg13g2_fill_2
X_3650_ _0491_ _0485_ _0453_ _0508_ VPWR VGND sg13g2_a21o_1
X_3581_ _0440_ _0432_ _0441_ VPWR VGND sg13g2_nor2b_1
X_5320_ net515 VPWR _2104_ VGND _2098_ _2102_ sg13g2_o21ai_1
XFILLER_6_871 VPWR VGND sg13g2_fill_1
X_5251_ _2043_ _2038_ _2041_ VPWR VGND sg13g2_xnor2_1
X_4202_ _1030_ _1031_ _1033_ _1034_ VPWR VGND sg13g2_or3_1
X_5182_ _1950_ _1944_ _1952_ _1976_ VPWR VGND sg13g2_a21o_1
X_4133_ _0970_ _0957_ _0972_ VPWR VGND sg13g2_xor2_1
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
X_4064_ _0905_ _0904_ _0902_ VPWR VGND sg13g2_nand2b_1
X_3015_ _2612_ _2603_ _2610_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_959 VPWR VGND sg13g2_decap_8
X_4966_ net798 net795 net846 net845 _1766_ VPWR VGND sg13g2_and4_1
X_4897_ _1703_ _1693_ _1704_ VPWR VGND sg13g2_nor2b_1
X_3917_ _0762_ _0718_ _0761_ VPWR VGND sg13g2_xnor2_1
X_3848_ _0695_ net917 net968 VPWR VGND sg13g2_nand2_1
X_3779_ _0624_ VPWR _0629_ VGND _0625_ _0627_ sg13g2_o21ai_1
X_5518_ _2257_ mac2.sum_lvl3_ff\[23\] mac2.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
X_5449_ net361 _2201_ _0041_ VPWR VGND sg13g2_xor2_1
XFILLER_28_786 VPWR VGND sg13g2_fill_2
XFILLER_43_712 VPWR VGND sg13g2_fill_2
XFILLER_15_414 VPWR VGND sg13g2_fill_2
XFILLER_42_200 VPWR VGND sg13g2_fill_1
XFILLER_15_458 VPWR VGND sg13g2_fill_1
XFILLER_24_981 VPWR VGND sg13g2_decap_8
XFILLER_30_439 VPWR VGND sg13g2_fill_1
XFILLER_10_152 VPWR VGND sg13g2_fill_1
XFILLER_10_185 VPWR VGND sg13g2_decap_4
XFILLER_19_731 VPWR VGND sg13g2_fill_2
XFILLER_38_539 VPWR VGND sg13g2_decap_8
XFILLER_46_561 VPWR VGND sg13g2_decap_4
XFILLER_18_241 VPWR VGND sg13g2_fill_1
X_4820_ _1628_ _1607_ _1630_ VPWR VGND sg13g2_xor2_1
X_4751_ _1563_ _1532_ _1561_ VPWR VGND sg13g2_xnor2_1
X_3702_ _0557_ _0558_ _0559_ VPWR VGND sg13g2_nor2_1
XFILLER_30_962 VPWR VGND sg13g2_decap_8
X_4682_ _1495_ _1487_ _1493_ VPWR VGND sg13g2_xnor2_1
X_3633_ _0492_ _0485_ _0491_ VPWR VGND sg13g2_xnor2_1
X_6421_ net1027 VGND VPWR net3 DP_1.I_range.out_data\[4\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_6352_ net1092 VGND VPWR _0142_ mac2.products_ff\[13\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3564_ _0378_ VPWR _0425_ VGND _0317_ _0379_ sg13g2_o21ai_1
X_5303_ net416 _2088_ _0008_ VPWR VGND sg13g2_xor2_1
X_6283_ net1023 VGND VPWR net74 mac1.sum_lvl3_ff\[28\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3495_ _0357_ net929 net986 VPWR VGND sg13g2_nand2_1
X_5234_ _2027_ _2006_ _2026_ VPWR VGND sg13g2_xnor2_1
X_5165_ _1960_ _1915_ _1958_ VPWR VGND sg13g2_xnor2_1
X_4116_ VGND VPWR _0925_ _0950_ _0955_ _0951_ sg13g2_a21oi_1
XFILLER_29_528 VPWR VGND sg13g2_fill_1
X_5096_ _1892_ _1891_ _1822_ _1893_ VPWR VGND sg13g2_a21o_1
X_4047_ _0889_ _0883_ _0888_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_200 VPWR VGND sg13g2_fill_2
XFILLER_25_712 VPWR VGND sg13g2_decap_4
X_5998_ net1069 VGND VPWR _0113_ mac1.products_ff\[7\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_4949_ _1748_ _1747_ _1742_ _1750_ VPWR VGND sg13g2_a21o_1
XFILLER_21_962 VPWR VGND sg13g2_decap_8
XFILLER_3_159 VPWR VGND sg13g2_fill_2
XFILLER_0_899 VPWR VGND sg13g2_decap_8
XFILLER_43_586 VPWR VGND sg13g2_fill_2
XFILLER_8_966 VPWR VGND sg13g2_decap_8
XFILLER_48_1024 VPWR VGND sg13g2_decap_4
X_3280_ _2868_ _2864_ _2869_ VPWR VGND sg13g2_xor2_1
X_5921_ net272 _0171_ VPWR VGND sg13g2_buf_1
XFILLER_0_1004 VPWR VGND sg13g2_decap_8
X_5852_ _2425_ _2428_ _2424_ _2547_ VPWR VGND sg13g2_nand3_1
XFILLER_34_586 VPWR VGND sg13g2_fill_1
X_4803_ _1613_ _1587_ _1611_ VPWR VGND sg13g2_xnor2_1
X_5783_ _2490_ _2486_ net760 VPWR VGND sg13g2_nand2b_1
X_2995_ _2594_ net956 net898 _0064_ VPWR VGND sg13g2_and3_2
X_4734_ _1546_ net826 net875 VPWR VGND sg13g2_nand2_1
X_4665_ _1477_ _1478_ _1448_ _1479_ VPWR VGND sg13g2_nand3_1
X_3616_ _0475_ net990 net1005 VPWR VGND sg13g2_nand2_1
X_6404_ net1057 VGND VPWR net138 mac2.sum_lvl1_ff\[37\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_4596_ _1408_ _1409_ _1372_ _1412_ VPWR VGND sg13g2_nand3_1
X_3547_ _0408_ net1010 net938 net978 net933 VPWR VGND sg13g2_a22oi_1
X_6335_ net1018 VGND VPWR net325 mac1.total_sum\[12\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3478_ _0341_ _0338_ _0340_ VPWR VGND sg13g2_nand2_1
X_6266_ net1035 VGND VPWR net208 mac2.sum_lvl1_ff\[79\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5217_ _2010_ _2009_ _2007_ VPWR VGND sg13g2_nand2b_1
X_6197_ net1064 VGND VPWR net131 mac1.sum_lvl2_ff\[21\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_5148_ _1907_ VPWR _1943_ VGND _1904_ _1908_ sg13g2_o21ai_1
X_5079_ net797 net794 net839 net997 _1876_ VPWR VGND sg13g2_and4_1
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_29_881 VPWR VGND sg13g2_decap_8
XFILLER_16_586 VPWR VGND sg13g2_fill_2
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
XFILLER_12_792 VPWR VGND sg13g2_fill_1
XFILLER_11_280 VPWR VGND sg13g2_fill_2
X_4450_ _1245_ VPWR _1275_ VGND _1243_ _1246_ sg13g2_o21ai_1
Xhold207 mac1.products_ff\[78\] VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold218 mac2.products_ff\[150\] VPWR VGND net258 sg13g2_dlygate4sd3_1
X_3401_ _2968_ _2981_ _2982_ VPWR VGND sg13g2_nor2b_1
Xhold229 DP_1.matrix\[80\] VPWR VGND net269 sg13g2_dlygate4sd3_1
X_4381_ _1208_ net868 net995 VPWR VGND sg13g2_nand2_1
X_6120_ net1092 VGND VPWR _0233_ DP_3.matrix\[41\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3332_ _2919_ _2918_ _2915_ VPWR VGND sg13g2_nand2b_1
X_3263_ _2852_ _2849_ _0095_ VPWR VGND sg13g2_xor2_1
X_6051_ net1085 VGND VPWR _0187_ DP_1.matrix\[43\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_3194_ _2785_ _2735_ _2783_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_100 VPWR VGND sg13g2_fill_2
X_5002_ _1797_ _1798_ _1800_ _1801_ VPWR VGND sg13g2_or3_1
X_5904_ _2579_ VPWR _0248_ VGND net761 _2580_ sg13g2_o21ai_1
XFILLER_35_873 VPWR VGND sg13g2_decap_8
X_5835_ net985 net753 _2536_ VPWR VGND sg13g2_nor2_1
XFILLER_14_16 VPWR VGND sg13g2_fill_2
X_5766_ _2473_ net271 net766 VPWR VGND sg13g2_nand2_1
X_5697_ _2406_ net771 _2405_ net764 net270 VPWR VGND sg13g2_a22oi_1
X_4717_ _1484_ _1529_ _1483_ _1530_ VPWR VGND sg13g2_nand3_1
X_4648_ _1431_ VPWR _1462_ VGND _1429_ _1432_ sg13g2_o21ai_1
X_4579_ _1393_ _1390_ _1395_ VPWR VGND sg13g2_xor2_1
X_6318_ net1029 VGND VPWR net56 mac2.sum_lvl3_ff\[31\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6249_ net1014 VGND VPWR net144 mac1.sum_lvl1_ff\[78\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_26_873 VPWR VGND sg13g2_decap_8
XFILLER_38_1012 VPWR VGND sg13g2_decap_8
XFILLER_41_821 VPWR VGND sg13g2_fill_2
XFILLER_9_538 VPWR VGND sg13g2_fill_2
XFILLER_5_788 VPWR VGND sg13g2_fill_2
XFILLER_1_983 VPWR VGND sg13g2_decap_8
XFILLER_49_954 VPWR VGND sg13g2_decap_8
XFILLER_36_626 VPWR VGND sg13g2_fill_1
Xhold90 mac2.sum_lvl1_ff\[49\] VPWR VGND net130 sg13g2_dlygate4sd3_1
X_3950_ _0793_ _0794_ _0795_ VPWR VGND sg13g2_and2_1
XFILLER_32_821 VPWR VGND sg13g2_fill_1
X_3881_ _0727_ _0723_ _0726_ VPWR VGND sg13g2_xnor2_1
X_5620_ mac2.total_sum\[10\] mac1.total_sum\[10\] _2336_ VPWR VGND sg13g2_xor2_1
X_5551_ _2278_ _2282_ _2283_ VPWR VGND sg13g2_nor2_1
X_4502_ _1309_ _1301_ _1308_ _1325_ VPWR VGND sg13g2_a21o_1
X_5482_ mac2.sum_lvl2_ff\[30\] mac2.sum_lvl2_ff\[11\] _2229_ VPWR VGND sg13g2_and2_1
X_4433_ _1257_ _1249_ _1259_ VPWR VGND sg13g2_xor2_1
X_4364_ _1192_ _1177_ _1191_ VPWR VGND sg13g2_nand2_1
X_6103_ net1064 VGND VPWR net57 mac1.sum_lvl1_ff\[2\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3315_ _2903_ _2882_ _2902_ VPWR VGND sg13g2_xnor2_1
X_4295_ _1123_ _1084_ _1124_ VPWR VGND sg13g2_xor2_1
X_6034_ net1037 VGND VPWR _0171_ DP_4.matrix\[80\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3246_ _2832_ _2834_ _2835_ _2836_ VPWR VGND sg13g2_nor3_1
XFILLER_6_1010 VPWR VGND sg13g2_decap_8
X_3177_ _2767_ _2766_ _2732_ _2769_ VPWR VGND sg13g2_a21o_1
XFILLER_27_659 VPWR VGND sg13g2_fill_1
XFILLER_41_128 VPWR VGND sg13g2_fill_1
XFILLER_34_191 VPWR VGND sg13g2_fill_1
X_5818_ _2524_ _2521_ _2523_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_898 VPWR VGND sg13g2_decap_4
X_5749_ net862 net779 _2456_ VPWR VGND sg13g2_nor2_1
XFILLER_46_924 VPWR VGND sg13g2_decap_8
XFILLER_18_637 VPWR VGND sg13g2_fill_1
XFILLER_18_659 VPWR VGND sg13g2_decap_8
XFILLER_14_810 VPWR VGND sg13g2_fill_2
XFILLER_14_854 VPWR VGND sg13g2_fill_2
XFILLER_41_695 VPWR VGND sg13g2_fill_1
X_3100_ _2693_ _2692_ _0101_ VPWR VGND sg13g2_xor2_1
XFILLER_1_791 VPWR VGND sg13g2_decap_8
X_4080_ _0920_ _0919_ _0921_ VPWR VGND sg13g2_nor2b_1
X_3031_ _2625_ _2626_ _2620_ _2627_ VPWR VGND sg13g2_nand3_1
XFILLER_37_902 VPWR VGND sg13g2_decap_8
XFILLER_37_979 VPWR VGND sg13g2_decap_8
X_4982_ _1754_ VPWR _1782_ VGND _1778_ _1779_ sg13g2_o21ai_1
X_3933_ _0778_ _0771_ _0776_ _0777_ VPWR VGND sg13g2_and3_1
X_3864_ _0711_ _0682_ _0710_ VPWR VGND sg13g2_nand2b_1
X_5603_ _2318_ _2321_ _2322_ _2323_ VPWR VGND sg13g2_nor3_1
X_3795_ _0644_ net970 net923 net971 net921 VPWR VGND sg13g2_a22oi_1
X_5534_ _2268_ net459 _0060_ VPWR VGND sg13g2_nor2b_1
X_5465_ mac2.sum_lvl2_ff\[7\] mac2.sum_lvl2_ff\[26\] _2216_ VPWR VGND sg13g2_xor2_1
XFILLER_28_1000 VPWR VGND sg13g2_decap_8
X_4416_ _1225_ _1218_ _1186_ _1242_ VPWR VGND sg13g2_a21o_1
X_5396_ _2155_ _2158_ net519 _2163_ VPWR VGND sg13g2_or3_1
X_4347_ _1174_ _1166_ _1175_ VPWR VGND sg13g2_nor2b_1
X_4278_ _1105_ _1106_ _1089_ _1108_ VPWR VGND sg13g2_nand3_1
X_3229_ _2784_ VPWR _2819_ VGND _2781_ _2785_ sg13g2_o21ai_1
X_6017_ net1086 VGND VPWR _0117_ mac1.products_ff\[78\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_28_902 VPWR VGND sg13g2_decap_8
XFILLER_43_927 VPWR VGND sg13g2_decap_8
XFILLER_27_456 VPWR VGND sg13g2_fill_1
XFILLER_28_979 VPWR VGND sg13g2_decap_8
XFILLER_42_437 VPWR VGND sg13g2_fill_2
XFILLER_36_990 VPWR VGND sg13g2_decap_8
Xheichips25_SDR_36 VPWR VGND uio_oe[3] sg13g2_tiehi
Xhold390 _0023_ VPWR VGND net430 sg13g2_dlygate4sd3_1
XFILLER_42_1008 VPWR VGND sg13g2_decap_8
Xfanout870 DP_3.matrix\[37\] net870 VPWR VGND sg13g2_buf_2
Xfanout892 net893 net892 VPWR VGND sg13g2_buf_8
Xfanout881 net493 net881 VPWR VGND sg13g2_buf_8
XFILLER_34_905 VPWR VGND sg13g2_decap_8
XFILLER_14_662 VPWR VGND sg13g2_decap_8
XFILLER_13_183 VPWR VGND sg13g2_fill_2
XFILLER_41_470 VPWR VGND sg13g2_fill_2
X_3580_ _0440_ _0433_ _0439_ VPWR VGND sg13g2_xnor2_1
X_5250_ _2042_ _2041_ _2038_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_371 VPWR VGND sg13g2_fill_1
X_4201_ _1033_ net862 net818 net863 net816 VPWR VGND sg13g2_a22oi_1
X_5181_ _1975_ _1972_ _0150_ VPWR VGND sg13g2_xor2_1
X_4132_ _0957_ _0970_ _0971_ VPWR VGND sg13g2_nor2_1
X_4063_ VGND VPWR _0904_ _0903_ _0853_ sg13g2_or2_1
X_3014_ _2611_ _2610_ _2603_ VPWR VGND sg13g2_nand2b_1
XFILLER_18_990 VPWR VGND sg13g2_decap_8
X_4965_ _1765_ net791 net849 VPWR VGND sg13g2_nand2_1
X_3916_ _0761_ _0753_ _0759_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_993 VPWR VGND sg13g2_decap_8
X_4896_ _1703_ _1679_ _1702_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_621 VPWR VGND sg13g2_decap_4
X_3847_ _0665_ VPWR _0694_ VGND _0663_ _0666_ sg13g2_o21ai_1
XFILLER_20_654 VPWR VGND sg13g2_fill_1
X_3778_ _0624_ _0625_ _0627_ _0628_ VPWR VGND sg13g2_nor3_1
X_5517_ VGND VPWR _2253_ _2255_ _2256_ _2254_ sg13g2_a21oi_1
X_6497_ net1031 VGND VPWR net16 DP_3.I_range.out_data\[6\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5448_ _2203_ mac2.sum_lvl2_ff\[22\] net360 VPWR VGND sg13g2_xnor2_1
X_5379_ _2147_ VPWR _2149_ VGND _2146_ _2148_ sg13g2_o21ai_1
XFILLER_16_949 VPWR VGND sg13g2_decap_8
XFILLER_43_746 VPWR VGND sg13g2_fill_1
XFILLER_24_960 VPWR VGND sg13g2_decap_8
XFILLER_30_429 VPWR VGND sg13g2_fill_2
XFILLER_11_643 VPWR VGND sg13g2_fill_2
XFILLER_3_886 VPWR VGND sg13g2_fill_1
XFILLER_34_735 VPWR VGND sg13g2_decap_4
XFILLER_33_234 VPWR VGND sg13g2_fill_2
XFILLER_30_941 VPWR VGND sg13g2_decap_8
X_4750_ _1562_ _1532_ _1561_ VPWR VGND sg13g2_nand2_1
X_3701_ VGND VPWR _0507_ _0528_ _0558_ _0530_ sg13g2_a21oi_1
X_4681_ _1494_ _1487_ _1493_ VPWR VGND sg13g2_nand2_1
X_3632_ _0490_ _0486_ _0491_ VPWR VGND sg13g2_xor2_1
X_6420_ net1027 VGND VPWR net2 DP_1.I_range.out_data\[3\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_6351_ net1092 VGND VPWR _0141_ mac2.products_ff\[12\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_5302_ net415 mac1.sum_lvl2_ff\[21\] _2090_ VPWR VGND sg13g2_xor2_1
X_3563_ _0421_ _0422_ _0352_ _0424_ VPWR VGND sg13g2_nand3_1
X_6282_ net1022 VGND VPWR net143 mac1.sum_lvl3_ff\[27\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3494_ _0356_ net986 net928 VPWR VGND sg13g2_nand2_1
X_5233_ _2026_ _2023_ _2024_ VPWR VGND sg13g2_xnor2_1
X_5164_ VGND VPWR _1959_ _1957_ _1916_ sg13g2_or2_1
X_4115_ _0926_ _0952_ _0954_ VPWR VGND sg13g2_and2_1
X_5095_ _1890_ _1889_ _1855_ _1892_ VPWR VGND sg13g2_a21o_1
X_4046_ _0887_ _0884_ _0888_ VPWR VGND sg13g2_xor2_1
X_5997_ net1067 VGND VPWR _0112_ mac1.products_ff\[6\] clknet_leaf_52_clk sg13g2_dfrbpq_1
XFILLER_21_941 VPWR VGND sg13g2_decap_8
X_4948_ _1747_ _1748_ _1742_ _1749_ VPWR VGND sg13g2_nand3_1
X_4879_ _1685_ _1686_ _1687_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_1018 VPWR VGND sg13g2_decap_8
XFILLER_48_849 VPWR VGND sg13g2_decap_8
XFILLER_43_510 VPWR VGND sg13g2_fill_1
XFILLER_43_543 VPWR VGND sg13g2_decap_4
XFILLER_43_532 VPWR VGND sg13g2_fill_2
XFILLER_15_267 VPWR VGND sg13g2_decap_4
XFILLER_8_945 VPWR VGND sg13g2_decap_8
XFILLER_7_433 VPWR VGND sg13g2_fill_1
XFILLER_11_462 VPWR VGND sg13g2_fill_2
XFILLER_12_985 VPWR VGND sg13g2_decap_8
XFILLER_48_1003 VPWR VGND sg13g2_decap_8
XFILLER_38_337 VPWR VGND sg13g2_fill_1
XFILLER_19_540 VPWR VGND sg13g2_decap_4
X_5920_ net273 _0170_ VPWR VGND sg13g2_buf_1
XFILLER_0_74 VPWR VGND sg13g2_fill_2
X_5851_ net930 net753 _2546_ VPWR VGND sg13g2_nor2_1
X_4802_ VGND VPWR _1612_ _1611_ _1587_ sg13g2_or2_1
X_5782_ VGND VPWR net1001 net760 _2489_ _2488_ sg13g2_a21oi_1
X_2994_ net958 net903 _0064_ VPWR VGND sg13g2_and2_1
X_4733_ _1545_ net879 net822 VPWR VGND sg13g2_nand2_1
XFILLER_9_83 VPWR VGND sg13g2_fill_2
X_6403_ net1057 VGND VPWR net163 mac2.sum_lvl1_ff\[36\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_4664_ _1455_ VPWR _1478_ VGND _1474_ _1476_ sg13g2_o21ai_1
X_3615_ _0447_ VPWR _0474_ VGND _0444_ _0448_ sg13g2_o21ai_1
X_4595_ _1411_ _1372_ _1408_ _1409_ VPWR VGND sg13g2_and3_1
X_3546_ net934 net978 net938 _0407_ VPWR VGND net1010 sg13g2_nand4_1
X_6334_ net1017 VGND VPWR net395 mac1.total_sum\[11\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_6265_ net1036 VGND VPWR net245 mac2.sum_lvl1_ff\[78\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5216_ VGND VPWR _2009_ _2008_ _1957_ sg13g2_or2_1
X_3477_ _0337_ _0336_ _0319_ _0340_ VPWR VGND sg13g2_a21o_1
X_6196_ net1045 VGND VPWR net96 mac1.sum_lvl2_ff\[20\] clknet_leaf_55_clk sg13g2_dfrbpq_1
XFILLER_28_48 VPWR VGND sg13g2_fill_1
XFILLER_29_304 VPWR VGND sg13g2_fill_2
XFILLER_29_326 VPWR VGND sg13g2_fill_1
X_5147_ _1929_ VPWR _1942_ VGND _1912_ _1930_ sg13g2_o21ai_1
X_5078_ _1875_ net791 net842 VPWR VGND sg13g2_nand2_1
X_4029_ _0872_ _0870_ _0871_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_893 VPWR VGND sg13g2_decap_8
XFILLER_37_392 VPWR VGND sg13g2_fill_1
XFILLER_5_937 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_fill_2
XFILLER_47_101 VPWR VGND sg13g2_fill_2
XFILLER_29_860 VPWR VGND sg13g2_decap_8
XFILLER_43_340 VPWR VGND sg13g2_fill_2
XFILLER_34_80 VPWR VGND sg13g2_fill_1
XFILLER_31_579 VPWR VGND sg13g2_fill_1
XFILLER_7_241 VPWR VGND sg13g2_fill_2
XFILLER_8_775 VPWR VGND sg13g2_fill_1
XFILLER_7_263 VPWR VGND sg13g2_fill_1
Xhold208 mac2.products_ff\[7\] VPWR VGND net248 sg13g2_dlygate4sd3_1
X_3400_ _2981_ _2969_ _2979_ VPWR VGND sg13g2_xnor2_1
Xhold219 mac1.products_ff\[145\] VPWR VGND net259 sg13g2_dlygate4sd3_1
X_4380_ _1180_ VPWR _1207_ VGND _1178_ _1181_ sg13g2_o21ai_1
X_3331_ _2917_ _2890_ _2918_ VPWR VGND sg13g2_xor2_1
X_3262_ _2852_ _2850_ _2851_ VPWR VGND sg13g2_nand2b_1
X_6050_ net1085 VGND VPWR _0186_ DP_1.matrix\[42\] clknet_leaf_48_clk sg13g2_dfrbpq_2
X_5001_ _1800_ net841 net797 net845 net793 VPWR VGND sg13g2_a22oi_1
X_3193_ VGND VPWR _2784_ _2782_ _2736_ sg13g2_or2_1
XFILLER_35_830 VPWR VGND sg13g2_fill_2
X_5903_ _2514_ _2510_ _2580_ VPWR VGND sg13g2_xor2_1
X_5834_ VGND VPWR net753 _2535_ _0175_ _2534_ sg13g2_a21oi_1
XFILLER_22_502 VPWR VGND sg13g2_decap_4
XFILLER_22_513 VPWR VGND sg13g2_fill_2
XFILLER_22_557 VPWR VGND sg13g2_fill_1
X_5765_ _2472_ _2471_ _2460_ VPWR VGND sg13g2_nand2b_1
X_5696_ net979 net962 net776 _2405_ VPWR VGND sg13g2_mux2_1
X_4716_ _1527_ _1528_ _1529_ VPWR VGND sg13g2_and2_1
X_4647_ _1461_ _1457_ _1460_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_929 VPWR VGND sg13g2_decap_8
X_6317_ net1028 VGND VPWR net85 mac2.sum_lvl3_ff\[30\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_4578_ _1394_ _1393_ _1390_ VPWR VGND sg13g2_nand2b_1
X_3529_ _0389_ _0349_ _0390_ VPWR VGND sg13g2_xor2_1
X_6248_ net1014 VGND VPWR net175 mac1.sum_lvl1_ff\[77\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_6179_ net1044 VGND VPWR net146 mac1.sum_lvl2_ff\[0\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_26_852 VPWR VGND sg13g2_decap_8
XFILLER_41_899 VPWR VGND sg13g2_decap_8
XFILLER_5_767 VPWR VGND sg13g2_fill_1
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_962 VPWR VGND sg13g2_decap_8
XFILLER_49_933 VPWR VGND sg13g2_decap_8
XFILLER_0_472 VPWR VGND sg13g2_fill_1
Xhold91 mac1.sum_lvl1_ff\[38\] VPWR VGND net131 sg13g2_dlygate4sd3_1
Xhold80 mac1.sum_lvl2_ff\[43\] VPWR VGND net120 sg13g2_dlygate4sd3_1
X_3880_ _0726_ _0689_ _0724_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_899 VPWR VGND sg13g2_decap_8
X_5550_ VPWR VGND net338 _2275_ mac2.sum_lvl3_ff\[29\] mac2.sum_lvl3_ff\[28\] _2282_
+ mac2.sum_lvl3_ff\[8\] sg13g2_a221oi_1
X_4501_ _1313_ _1315_ _1324_ VPWR VGND sg13g2_and2_1
XFILLER_8_550 VPWR VGND sg13g2_fill_2
X_5481_ _2228_ net545 _0033_ VPWR VGND sg13g2_xor2_1
X_4432_ _1257_ _1249_ _1258_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_594 VPWR VGND sg13g2_fill_1
X_4363_ _1190_ _1183_ _1191_ VPWR VGND sg13g2_xor2_1
X_3314_ _2902_ _2899_ _2900_ VPWR VGND sg13g2_xnor2_1
X_6102_ net1055 VGND VPWR _0221_ DP_3.matrix\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4294_ _1123_ net868 net803 VPWR VGND sg13g2_nand2_1
X_6033_ net1092 VGND VPWR _0170_ DP_4.matrix\[44\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3245_ _2835_ net941 net895 net945 net893 VPWR VGND sg13g2_a22oi_1
X_3176_ _2766_ _2767_ _2732_ _2768_ VPWR VGND sg13g2_nand3_1
XFILLER_23_833 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_61_clk clknet_4_8_0_clk clknet_leaf_61_clk VPWR VGND sg13g2_buf_8
X_5817_ _2523_ _2522_ net768 net766 net782 VPWR VGND sg13g2_a22oi_1
X_5748_ _2455_ net274 net765 VPWR VGND sg13g2_nand2_1
X_5679_ _2388_ _2386_ _2387_ _2385_ net770 VPWR VGND sg13g2_a22oi_1
XFILLER_46_903 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_52_clk clknet_4_8_0_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
XFILLER_40_151 VPWR VGND sg13g2_decap_8
XFILLER_41_674 VPWR VGND sg13g2_fill_1
XFILLER_13_387 VPWR VGND sg13g2_fill_1
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_785 VPWR VGND sg13g2_decap_8
X_3030_ _2621_ VPWR _2626_ VGND _2622_ _2624_ sg13g2_o21ai_1
XFILLER_49_796 VPWR VGND sg13g2_fill_2
XFILLER_37_958 VPWR VGND sg13g2_decap_8
X_4981_ _1754_ _1778_ _1779_ _1781_ VPWR VGND sg13g2_nor3_1
X_3932_ _0772_ VPWR _0777_ VGND _0773_ _0775_ sg13g2_o21ai_1
XFILLER_16_181 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_43_clk clknet_4_11_0_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_3863_ _0710_ _0686_ _0709_ VPWR VGND sg13g2_xnor2_1
X_5602_ VPWR VGND _2316_ _2315_ _2314_ mac1.total_sum\[5\] _2322_ mac2.total_sum\[5\]
+ sg13g2_a221oi_1
XFILLER_20_858 VPWR VGND sg13g2_fill_1
X_3794_ net921 net971 net923 _0643_ VPWR VGND net970 sg13g2_nand4_1
X_5533_ net458 VPWR _2269_ VGND _2263_ _2267_ sg13g2_o21ai_1
X_5464_ _2215_ mac2.sum_lvl2_ff\[26\] net506 VPWR VGND sg13g2_nand2_1
X_5395_ net519 VPWR _2162_ VGND _2155_ _2158_ sg13g2_o21ai_1
X_4415_ _1227_ VPWR _1241_ VGND _1216_ _1228_ sg13g2_o21ai_1
X_4346_ _1174_ _1167_ _1173_ VPWR VGND sg13g2_xnor2_1
X_4277_ _1107_ _1089_ _1105_ _1106_ VPWR VGND sg13g2_and3_1
X_6016_ net1078 VGND VPWR _0126_ mac1.products_ff\[77\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_3228_ _2805_ VPWR _2818_ VGND _2789_ _2806_ sg13g2_o21ai_1
XFILLER_39_251 VPWR VGND sg13g2_fill_1
X_3159_ _2711_ VPWR _2751_ VGND _2709_ _2712_ sg13g2_o21ai_1
XFILLER_28_958 VPWR VGND sg13g2_decap_8
XFILLER_43_906 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_34_clk clknet_4_15_0_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_23_685 VPWR VGND sg13g2_fill_1
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_324 VPWR VGND sg13g2_fill_2
Xheichips25_SDR_37 VPWR VGND uio_oe[4] sg13g2_tiehi
Xhold380 _0059_ VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold391 DP_2.matrix\[4\] VPWR VGND net431 sg13g2_dlygate4sd3_1
Xfanout860 net472 net860 VPWR VGND sg13g2_buf_8
Xfanout893 net307 net893 VPWR VGND sg13g2_buf_8
Xfanout871 net363 net871 VPWR VGND sg13g2_buf_8
Xfanout882 net883 net882 VPWR VGND sg13g2_buf_8
XFILLER_45_221 VPWR VGND sg13g2_fill_1
XFILLER_27_980 VPWR VGND sg13g2_decap_8
XFILLER_33_416 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_25_clk clknet_4_7_0_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_33_438 VPWR VGND sg13g2_fill_1
XFILLER_42_994 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_fill_1
XFILLER_47_4 VPWR VGND sg13g2_fill_2
X_4200_ net816 net863 net818 _1032_ VPWR VGND net862 sg13g2_nand4_1
X_5180_ _1975_ _1973_ _1974_ VPWR VGND sg13g2_nand2b_1
X_4131_ _0968_ _0958_ _0970_ VPWR VGND sg13g2_xor2_1
X_4062_ _0903_ net910 net1009 VPWR VGND sg13g2_nand2_1
XFILLER_49_593 VPWR VGND sg13g2_decap_8
X_3013_ _2608_ _2609_ _2610_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_416 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_16_clk clknet_4_4_0_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_4964_ _1745_ VPWR _1764_ VGND _1743_ _1746_ sg13g2_o21ai_1
X_3915_ _0760_ _0753_ _0759_ VPWR VGND sg13g2_nand2_1
XFILLER_33_972 VPWR VGND sg13g2_decap_8
X_4895_ _1700_ _1699_ _1702_ VPWR VGND sg13g2_xor2_1
XFILLER_32_482 VPWR VGND sg13g2_fill_2
X_3846_ _0693_ _0688_ _0691_ VPWR VGND sg13g2_xnor2_1
X_3777_ _0627_ net972 net924 net973 net918 VPWR VGND sg13g2_a22oi_1
X_6496_ net1031 VGND VPWR DP_3.I_range.data_plus_4\[6\] DP_3.I_range.out_data\[5\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5516_ net452 _2253_ _0056_ VPWR VGND sg13g2_xor2_1
X_5447_ _2202_ mac2.sum_lvl2_ff\[22\] net360 VPWR VGND sg13g2_nand2_1
X_5378_ net384 _2146_ _0025_ VPWR VGND sg13g2_xor2_1
X_4329_ _1155_ _1156_ _1087_ _1158_ VPWR VGND sg13g2_nand3_1
XFILLER_28_744 VPWR VGND sg13g2_fill_2
XFILLER_43_714 VPWR VGND sg13g2_fill_1
XFILLER_28_788 VPWR VGND sg13g2_fill_1
XFILLER_10_110 VPWR VGND sg13g2_fill_1
XFILLER_23_471 VPWR VGND sg13g2_fill_2
XFILLER_19_733 VPWR VGND sg13g2_fill_1
XFILLER_34_747 VPWR VGND sg13g2_fill_1
XFILLER_18_1011 VPWR VGND sg13g2_decap_8
XFILLER_42_791 VPWR VGND sg13g2_fill_1
XFILLER_15_994 VPWR VGND sg13g2_decap_8
X_3700_ _0557_ _0536_ _0556_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_920 VPWR VGND sg13g2_decap_8
X_4680_ _1493_ _1488_ _1491_ VPWR VGND sg13g2_xnor2_1
X_3631_ _0490_ _0445_ _0488_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_997 VPWR VGND sg13g2_decap_8
X_3562_ _0422_ _0421_ _0352_ _0423_ VPWR VGND sg13g2_a21o_1
X_6350_ net1090 VGND VPWR _0140_ mac2.products_ff\[11\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_5301_ mac1.sum_lvl2_ff\[21\] net415 _2089_ VPWR VGND sg13g2_and2_1
X_6281_ net1022 VGND VPWR net106 mac1.sum_lvl3_ff\[26\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3493_ _0355_ net990 net927 VPWR VGND sg13g2_nand2_1
X_5232_ _2024_ _2023_ _2025_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5163_ _1958_ net789 net838 VPWR VGND sg13g2_nand2_1
XFILLER_25_1015 VPWR VGND sg13g2_decap_8
X_4114_ _0953_ _0952_ _0120_ VPWR VGND sg13g2_xor2_1
X_5094_ _1889_ _1890_ _1855_ _1891_ VPWR VGND sg13g2_nand3_1
XFILLER_17_28 VPWR VGND sg13g2_fill_2
X_4045_ _0887_ _0842_ _0885_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_541 VPWR VGND sg13g2_decap_8
XFILLER_37_574 VPWR VGND sg13g2_fill_2
X_5996_ net1064 VGND VPWR _0105_ mac1.products_ff\[5\] clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_33_27 VPWR VGND sg13g2_fill_2
X_4947_ _1743_ VPWR _1748_ VGND _1744_ _1746_ sg13g2_o21ai_1
X_4878_ _1686_ _1667_ _1684_ VPWR VGND sg13g2_nand2_1
X_3829_ _0677_ _0638_ _0674_ _0675_ VPWR VGND sg13g2_and3_1
XFILLER_21_997 VPWR VGND sg13g2_decap_8
X_6479_ net1013 VGND VPWR net541 mac2.total_sum\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_12_964 VPWR VGND sg13g2_decap_8
XFILLER_7_489 VPWR VGND sg13g2_fill_1
XFILLER_7_478 VPWR VGND sg13g2_fill_2
XFILLER_2_161 VPWR VGND sg13g2_fill_2
XFILLER_48_90 VPWR VGND sg13g2_fill_1
XFILLER_47_883 VPWR VGND sg13g2_decap_8
XFILLER_34_533 VPWR VGND sg13g2_fill_2
X_5850_ VGND VPWR net754 _2545_ _0197_ _2544_ sg13g2_a21oi_1
X_5781_ _2451_ net760 _2488_ VPWR VGND sg13g2_nor2_1
X_2993_ VPWR _2593_ net995 VGND sg13g2_inv_1
X_4801_ _1611_ net826 net1002 VPWR VGND sg13g2_nand2_1
X_4732_ _1513_ VPWR _1544_ VGND _1504_ _1514_ sg13g2_o21ai_1
X_4663_ _1455_ _1474_ _1476_ _1477_ VPWR VGND sg13g2_or3_1
X_6402_ net1093 VGND VPWR net264 mac2.sum_lvl1_ff\[15\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3614_ _0437_ VPWR _0473_ VGND _0434_ _0438_ sg13g2_o21ai_1
X_4594_ VGND VPWR _1408_ _1409_ _1410_ _1372_ sg13g2_a21oi_1
X_3545_ net938 net933 net978 net1010 _0406_ VPWR VGND sg13g2_and4_1
X_6333_ net1017 VGND VPWR net379 mac1.total_sum\[10\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3476_ VGND VPWR _0336_ _0337_ _0339_ _0319_ sg13g2_a21oi_1
X_6264_ net1036 VGND VPWR net185 mac2.sum_lvl1_ff\[77\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5215_ _2008_ net785 net997 VPWR VGND sg13g2_nand2_1
X_6195_ net1043 VGND VPWR net197 mac1.sum_lvl2_ff\[19\] clknet_leaf_62_clk sg13g2_dfrbpq_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
X_5146_ _1909_ _1903_ _1911_ _1941_ VPWR VGND sg13g2_a21o_1
X_5077_ _1834_ VPWR _1874_ VGND _1832_ _1835_ sg13g2_o21ai_1
X_4028_ VGND VPWR _0793_ _0833_ _0871_ _0834_ sg13g2_a21oi_1
XFILLER_38_872 VPWR VGND sg13g2_decap_8
XFILLER_25_566 VPWR VGND sg13g2_fill_2
XFILLER_25_577 VPWR VGND sg13g2_decap_4
X_5979_ net796 _0261_ VPWR VGND sg13g2_buf_1
XFILLER_13_739 VPWR VGND sg13g2_fill_2
XFILLER_12_249 VPWR VGND sg13g2_fill_2
XFILLER_20_293 VPWR VGND sg13g2_decap_4
XFILLER_47_157 VPWR VGND sg13g2_fill_1
XFILLER_44_886 VPWR VGND sg13g2_decap_8
XFILLER_16_588 VPWR VGND sg13g2_fill_1
XFILLER_12_772 VPWR VGND sg13g2_fill_2
XFILLER_11_282 VPWR VGND sg13g2_fill_1
Xhold209 mac1.products_ff\[138\] VPWR VGND net249 sg13g2_dlygate4sd3_1
X_3330_ _2917_ net889 net943 VPWR VGND sg13g2_nand2_1
XFILLER_4_982 VPWR VGND sg13g2_decap_8
X_3261_ VGND VPWR _2773_ _2813_ _2851_ _2814_ sg13g2_a21oi_1
X_5000_ net793 net845 net797 _1799_ VPWR VGND net842 sg13g2_nand4_1
X_3192_ _2783_ net953 net889 VPWR VGND sg13g2_nand2_1
XFILLER_22_1018 VPWR VGND sg13g2_decap_8
XFILLER_38_157 VPWR VGND sg13g2_fill_2
X_5902_ _2579_ net824 net761 VPWR VGND sg13g2_nand2_1
X_5833_ _2394_ _2382_ _2535_ VPWR VGND sg13g2_xor2_1
XFILLER_14_18 VPWR VGND sg13g2_fill_1
XFILLER_22_525 VPWR VGND sg13g2_decap_8
X_5764_ _2470_ _2468_ _2471_ VPWR VGND sg13g2_nor2b_1
X_5695_ _2404_ _2401_ _2403_ VPWR VGND sg13g2_nand2b_1
X_4715_ _1525_ _1524_ _1526_ _1528_ VPWR VGND sg13g2_a21o_1
X_4646_ _1460_ _1423_ _1458_ VPWR VGND sg13g2_xnor2_1
X_4577_ _1392_ _1371_ _1393_ VPWR VGND sg13g2_xor2_1
XFILLER_2_908 VPWR VGND sg13g2_decap_8
X_6316_ net1028 VGND VPWR net113 mac2.sum_lvl3_ff\[29\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3528_ _0389_ net990 net926 VPWR VGND sg13g2_nand2_1
X_6247_ net1014 VGND VPWR net212 mac1.sum_lvl1_ff\[76\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3459_ _0322_ net988 net929 VPWR VGND sg13g2_nand2_1
X_6178_ net1083 VGND VPWR net60 mac1.sum_lvl1_ff\[51\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5129_ _1923_ _1924_ _1925_ VPWR VGND sg13g2_nor2_1
XFILLER_26_820 VPWR VGND sg13g2_decap_8
XFILLER_41_878 VPWR VGND sg13g2_decap_8
XFILLER_45_1007 VPWR VGND sg13g2_decap_8
XFILLER_1_941 VPWR VGND sg13g2_decap_8
XFILLER_49_912 VPWR VGND sg13g2_decap_8
XFILLER_49_989 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_fill_2
Xhold81 mac2.products_ff\[82\] VPWR VGND net121 sg13g2_dlygate4sd3_1
Xhold70 mac1.sum_lvl1_ff\[13\] VPWR VGND net110 sg13g2_dlygate4sd3_1
Xhold92 mac2.products_ff\[144\] VPWR VGND net132 sg13g2_dlygate4sd3_1
XFILLER_16_363 VPWR VGND sg13g2_fill_1
XFILLER_43_193 VPWR VGND sg13g2_fill_2
XFILLER_32_878 VPWR VGND sg13g2_decap_8
X_4500_ _1321_ _1297_ _1322_ _1323_ VPWR VGND sg13g2_a21o_1
X_5480_ _2223_ _2227_ _2228_ VPWR VGND sg13g2_nor2_1
X_4431_ _1257_ _1250_ _1256_ VPWR VGND sg13g2_xnor2_1
X_4362_ _1190_ _1184_ _1188_ VPWR VGND sg13g2_xnor2_1
X_3313_ _2900_ _2899_ _2901_ VPWR VGND sg13g2_nor2b_1
X_6101_ net1055 VGND VPWR _0220_ DP_3.matrix\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_4293_ _1122_ net868 net801 VPWR VGND sg13g2_nand2_1
X_6032_ net1075 VGND VPWR _0169_ DP_4.matrix\[8\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3244_ net895 net892 net945 net942 _2834_ VPWR VGND sg13g2_and4_1
XFILLER_20_0 VPWR VGND sg13g2_fill_2
XFILLER_39_433 VPWR VGND sg13g2_fill_1
X_3175_ _2742_ VPWR _2767_ VGND _2763_ _2765_ sg13g2_o21ai_1
Xfanout1090 net1091 net1090 VPWR VGND sg13g2_buf_8
XFILLER_34_160 VPWR VGND sg13g2_fill_1
XFILLER_41_119 VPWR VGND sg13g2_fill_1
X_5816_ net802 net820 net779 _2522_ VPWR VGND sg13g2_mux2_1
X_5747_ _2446_ net778 _2454_ VPWR VGND sg13g2_nor2_1
X_5678_ net770 VPWR _2387_ VGND net975 net774 sg13g2_o21ai_1
X_4629_ _1444_ _1420_ _1443_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_959 VPWR VGND sg13g2_decap_8
XFILLER_14_812 VPWR VGND sg13g2_fill_1
XFILLER_26_683 VPWR VGND sg13g2_decap_4
XFILLER_14_856 VPWR VGND sg13g2_fill_1
XFILLER_12_1006 VPWR VGND sg13g2_decap_8
XFILLER_49_764 VPWR VGND sg13g2_decap_8
XFILLER_37_937 VPWR VGND sg13g2_decap_8
XFILLER_36_469 VPWR VGND sg13g2_decap_4
X_4980_ _1776_ _1777_ _1740_ _1780_ VPWR VGND sg13g2_nand3_1
X_3931_ _0772_ _0773_ _0775_ _0776_ VPWR VGND sg13g2_or3_1
X_3862_ _0709_ _0706_ _0708_ VPWR VGND sg13g2_nand2_1
X_5601_ _2321_ mac1.total_sum\[6\] mac2.total_sum\[6\] VPWR VGND sg13g2_xnor2_1
XFILLER_31_185 VPWR VGND sg13g2_fill_2
XFILLER_32_697 VPWR VGND sg13g2_fill_2
XFILLER_9_860 VPWR VGND sg13g2_fill_2
X_3793_ net923 DP_2.matrix\[37\] net972 net970 _0642_ VPWR VGND sg13g2_and4_1
XFILLER_9_871 VPWR VGND sg13g2_fill_2
X_5532_ _2263_ net458 _2267_ _2268_ VPWR VGND sg13g2_nor3_1
XFILLER_9_893 VPWR VGND sg13g2_decap_4
X_5463_ _2213_ net526 _0044_ VPWR VGND sg13g2_nor2b_2
X_5394_ net518 mac1.sum_lvl3_ff\[27\] _2161_ VPWR VGND sg13g2_xor2_1
X_4414_ _1213_ _1207_ _1215_ _1240_ VPWR VGND sg13g2_a21o_1
X_4345_ _1172_ _1168_ _1173_ VPWR VGND sg13g2_xor2_1
X_4276_ _1094_ VPWR _1106_ VGND _1102_ _1104_ sg13g2_o21ai_1
X_3227_ _2786_ _2780_ _2788_ _2817_ VPWR VGND sg13g2_a21o_1
X_6015_ net1078 VGND VPWR _0125_ mac1.products_ff\[76\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3158_ _2750_ _2749_ _2748_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_937 VPWR VGND sg13g2_decap_8
X_3089_ _2680_ _2679_ _2674_ _2683_ VPWR VGND sg13g2_a21o_1
XFILLER_35_1006 VPWR VGND sg13g2_decap_8
Xheichips25_SDR_38 VPWR VGND uio_oe[5] sg13g2_tiehi
Xhold370 _2193_ VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold381 DP_3.matrix\[75\] VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold392 _2551_ VPWR VGND net432 sg13g2_dlygate4sd3_1
Xfanout861 net862 net861 VPWR VGND sg13g2_buf_8
Xfanout850 net851 net850 VPWR VGND sg13g2_buf_8
Xfanout872 DP_3.matrix\[7\] net872 VPWR VGND sg13g2_buf_8
Xfanout894 net895 net894 VPWR VGND sg13g2_buf_8
Xfanout883 net498 net883 VPWR VGND sg13g2_buf_8
XFILLER_19_959 VPWR VGND sg13g2_decap_8
XFILLER_42_973 VPWR VGND sg13g2_decap_8
XFILLER_13_152 VPWR VGND sg13g2_fill_1
XFILLER_13_185 VPWR VGND sg13g2_fill_1
XFILLER_41_472 VPWR VGND sg13g2_fill_1
XFILLER_41_494 VPWR VGND sg13g2_fill_1
XFILLER_13_196 VPWR VGND sg13g2_decap_4
XFILLER_42_92 VPWR VGND sg13g2_decap_8
X_4130_ _0968_ _0958_ _0969_ VPWR VGND sg13g2_nor2b_1
X_4061_ _0902_ net1009 net913 net961 net910 VPWR VGND sg13g2_a22oi_1
XFILLER_49_572 VPWR VGND sg13g2_fill_2
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
X_3012_ _2604_ VPWR _2609_ VGND _2605_ _2607_ sg13g2_o21ai_1
XFILLER_36_244 VPWR VGND sg13g2_fill_1
X_4963_ _1761_ _1758_ _1763_ VPWR VGND sg13g2_xor2_1
X_3914_ _0759_ _0754_ _0757_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_951 VPWR VGND sg13g2_decap_8
X_4894_ _1701_ _1699_ _1700_ VPWR VGND sg13g2_nand2_1
XFILLER_32_461 VPWR VGND sg13g2_fill_1
X_3845_ _0692_ _0691_ _0688_ VPWR VGND sg13g2_nand2b_1
X_3776_ net918 net973 net924 _0626_ VPWR VGND net972 sg13g2_nand4_1
X_6495_ net1031 VGND VPWR net15 DP_3.I_range.out_data\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5515_ net451 mac2.sum_lvl3_ff\[22\] _2255_ VPWR VGND sg13g2_xor2_1
X_5446_ VGND VPWR _2198_ net321 _2201_ _2199_ sg13g2_a21oi_1
X_5377_ _2148_ mac1.sum_lvl3_ff\[23\] net383 VPWR VGND sg13g2_xnor2_1
X_4328_ _1156_ _1155_ _1087_ _1157_ VPWR VGND sg13g2_a21o_1
X_4259_ _1070_ _1060_ _1068_ _1089_ VPWR VGND sg13g2_a21o_1
XFILLER_27_266 VPWR VGND sg13g2_decap_4
XFILLER_42_258 VPWR VGND sg13g2_fill_2
XFILLER_24_995 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_4
XFILLER_14_450 VPWR VGND sg13g2_fill_2
XFILLER_15_973 VPWR VGND sg13g2_decap_8
XFILLER_14_461 VPWR VGND sg13g2_fill_2
X_3630_ VGND VPWR _0489_ _0487_ _0446_ sg13g2_or2_1
XFILLER_30_976 VPWR VGND sg13g2_decap_8
X_3561_ _0420_ _0419_ _0385_ _0422_ VPWR VGND sg13g2_a21o_1
X_5300_ _2085_ VPWR _2088_ VGND _2084_ _2086_ sg13g2_o21ai_1
X_6280_ net1022 VGND VPWR net120 mac1.sum_lvl3_ff\[25\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3492_ _0335_ _0325_ _0333_ _0354_ VPWR VGND sg13g2_a21o_1
X_5231_ VGND VPWR _1978_ _1983_ _2024_ _1997_ sg13g2_a21oi_1
X_5162_ _1957_ net787 net838 VPWR VGND sg13g2_nand2_2
X_4113_ _0953_ _0925_ _0931_ VPWR VGND sg13g2_nand2_1
X_5093_ _1865_ VPWR _1890_ VGND _1886_ _1888_ sg13g2_o21ai_1
X_4044_ VGND VPWR _0886_ _0885_ _0842_ sg13g2_or2_1
XFILLER_37_586 VPWR VGND sg13g2_fill_2
X_5995_ net1064 VGND VPWR _0073_ mac1.products_ff\[4\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_4946_ _1743_ _1744_ _1746_ _1747_ VPWR VGND sg13g2_or3_1
X_4877_ _1667_ _1684_ _1685_ VPWR VGND sg13g2_nor2_1
X_3828_ VGND VPWR _0674_ _0675_ _0676_ _0638_ sg13g2_a21oi_1
XFILLER_21_976 VPWR VGND sg13g2_decap_8
XFILLER_20_486 VPWR VGND sg13g2_fill_2
X_3759_ _0613_ _0607_ _0612_ VPWR VGND sg13g2_xnor2_1
X_6478_ net1016 VGND VPWR net460 mac2.total_sum\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_5429_ mac1.sum_lvl3_ff\[34\] net373 _2189_ VPWR VGND sg13g2_nor2_1
XFILLER_28_520 VPWR VGND sg13g2_fill_2
XFILLER_43_501 VPWR VGND sg13g2_decap_8
XFILLER_43_534 VPWR VGND sg13g2_fill_1
XFILLER_12_943 VPWR VGND sg13g2_decap_8
XFILLER_11_464 VPWR VGND sg13g2_fill_1
XFILLER_11_497 VPWR VGND sg13g2_fill_2
XFILLER_0_1018 VPWR VGND sg13g2_decap_8
XFILLER_19_597 VPWR VGND sg13g2_fill_1
X_4800_ _1610_ DP_4.matrix\[5\] net875 VPWR VGND sg13g2_nand2_1
X_2992_ VPWR _2592_ net999 VGND sg13g2_inv_1
X_5780_ DP_3.Q_range.out_data\[3\] _2452_ _2587_ _2487_ VPWR VGND _2453_ sg13g2_nand4_1
X_4731_ _1541_ _1533_ _1543_ VPWR VGND sg13g2_xor2_1
XFILLER_9_85 VPWR VGND sg13g2_fill_1
X_4662_ VGND VPWR _1472_ _1473_ _1476_ _1456_ sg13g2_a21oi_1
X_6401_ net1093 VGND VPWR net262 mac2.sum_lvl1_ff\[14\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3613_ _0459_ VPWR _0472_ VGND _0442_ _0460_ sg13g2_o21ai_1
X_4593_ _1407_ _1406_ _1389_ _1409_ VPWR VGND sg13g2_a21o_1
X_3544_ _0405_ net930 net981 VPWR VGND sg13g2_nand2_1
X_6332_ net1017 VGND VPWR net295 mac1.total_sum\[9\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3475_ _0336_ _0337_ _0319_ _0338_ VPWR VGND sg13g2_nand3_1
X_6263_ net1050 VGND VPWR net255 mac2.sum_lvl1_ff\[76\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5214_ _2007_ net997 net787 net838 net786 VPWR VGND sg13g2_a22oi_1
X_6194_ net1096 VGND VPWR net100 mac1.sum_lvl2_ff\[15\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5145_ _1940_ _1939_ _0159_ VPWR VGND sg13g2_xor2_1
X_5076_ _1873_ _1867_ _1872_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_309 VPWR VGND sg13g2_fill_2
X_4027_ _0750_ _0795_ _0749_ _0870_ VPWR VGND _0835_ sg13g2_nand4_1
XFILLER_44_49 VPWR VGND sg13g2_fill_1
X_5978_ net800 _0260_ VPWR VGND sg13g2_buf_1
XFILLER_40_504 VPWR VGND sg13g2_decap_8
X_4929_ _1726_ VPWR _1731_ VGND _1727_ _1729_ sg13g2_o21ai_1
XFILLER_47_103 VPWR VGND sg13g2_fill_1
XFILLER_47_114 VPWR VGND sg13g2_fill_1
XFILLER_29_895 VPWR VGND sg13g2_decap_8
XFILLER_31_537 VPWR VGND sg13g2_fill_1
XFILLER_8_722 VPWR VGND sg13g2_fill_1
XFILLER_8_711 VPWR VGND sg13g2_fill_2
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_766 VPWR VGND sg13g2_fill_2
XFILLER_7_243 VPWR VGND sg13g2_fill_1
XFILLER_7_287 VPWR VGND sg13g2_fill_1
XFILLER_4_961 VPWR VGND sg13g2_decap_8
X_3260_ _2730_ _2775_ _2729_ _2850_ VPWR VGND _2815_ sg13g2_nand4_1
X_3191_ _2782_ net953 net887 VPWR VGND sg13g2_nand2_1
X_5901_ _2578_ VPWR _0247_ VGND net762 _2577_ sg13g2_o21ai_1
X_5832_ net987 net753 _2534_ VPWR VGND sg13g2_nor2_1
XFILLER_34_364 VPWR VGND sg13g2_fill_2
XFILLER_35_887 VPWR VGND sg13g2_decap_8
XFILLER_34_397 VPWR VGND sg13g2_fill_2
X_5763_ _2470_ _2469_ net767 net765 net851 VPWR VGND sg13g2_a22oi_1
X_4714_ _1525_ _1526_ _1524_ _1527_ VPWR VGND sg13g2_nand3_1
X_5694_ _2403_ net771 _2402_ net764 net278 VPWR VGND sg13g2_a22oi_1
X_4645_ VGND VPWR _1459_ _1458_ _1423_ sg13g2_or2_1
X_4576_ _1392_ net882 net825 VPWR VGND sg13g2_nand2_1
X_3527_ _0388_ net990 net925 VPWR VGND sg13g2_nand2_1
X_6315_ net1020 VGND VPWR net137 mac2.sum_lvl3_ff\[28\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6246_ net1024 VGND VPWR net161 mac1.sum_lvl1_ff\[75\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_3458_ _0321_ net988 net928 VPWR VGND sg13g2_nand2_1
XFILLER_39_38 VPWR VGND sg13g2_decap_4
X_3389_ VGND VPWR _2963_ _2966_ _2970_ _2964_ sg13g2_a21oi_1
X_6177_ net1084 VGND VPWR net75 mac1.sum_lvl1_ff\[50\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5128_ _1924_ net998 net793 net838 net791 VPWR VGND sg13g2_a22oi_1
XFILLER_44_117 VPWR VGND sg13g2_fill_1
X_5059_ _1828_ VPWR _1856_ VGND _1825_ _1829_ sg13g2_o21ai_1
XFILLER_26_887 VPWR VGND sg13g2_decap_8
XFILLER_38_1026 VPWR VGND sg13g2_fill_2
XFILLER_1_920 VPWR VGND sg13g2_decap_8
XFILLER_1_997 VPWR VGND sg13g2_decap_8
XFILLER_49_968 VPWR VGND sg13g2_decap_8
Xhold60 mac1.sum_lvl1_ff\[15\] VPWR VGND net100 sg13g2_dlygate4sd3_1
Xhold71 mac2.products_ff\[8\] VPWR VGND net111 sg13g2_dlygate4sd3_1
Xhold82 mac2.products_ff\[5\] VPWR VGND net122 sg13g2_dlygate4sd3_1
Xhold93 mac2.sum_lvl1_ff\[2\] VPWR VGND net133 sg13g2_dlygate4sd3_1
XFILLER_28_180 VPWR VGND sg13g2_decap_8
XFILLER_45_92 VPWR VGND sg13g2_fill_2
XFILLER_44_684 VPWR VGND sg13g2_fill_1
XFILLER_16_353 VPWR VGND sg13g2_fill_2
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_8_552 VPWR VGND sg13g2_fill_1
X_4430_ _1255_ _1251_ _1256_ VPWR VGND sg13g2_xor2_1
X_6100_ net1045 VGND VPWR net198 mac1.sum_lvl1_ff\[1\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_4361_ _1189_ _1184_ _1188_ VPWR VGND sg13g2_nand2_1
XFILLER_4_791 VPWR VGND sg13g2_fill_1
X_3312_ VGND VPWR _2855_ _2860_ _2900_ _2873_ sg13g2_a21oi_1
X_4292_ _1121_ net871 net995 VPWR VGND sg13g2_nand2_1
X_6031_ net1037 VGND VPWR _0168_ DP_3.matrix\[80\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3243_ _2833_ net893 net943 VPWR VGND sg13g2_nand2_1
XFILLER_6_1024 VPWR VGND sg13g2_decap_4
X_3174_ _2742_ _2763_ _2765_ _2766_ VPWR VGND sg13g2_or3_1
Xfanout1080 net1082 net1080 VPWR VGND sg13g2_buf_8
Xfanout1091 net1097 net1091 VPWR VGND sg13g2_buf_8
XFILLER_23_813 VPWR VGND sg13g2_fill_2
X_5815_ _2516_ _2520_ _2521_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_835 VPWR VGND sg13g2_fill_1
X_5746_ DP_3.I_range.out_data\[6\] DP_3.I_range.out_data\[2\] _2588_ DP_3.I_range.out_data\[4\]
+ _2453_ VPWR VGND sg13g2_nor4_1
XFILLER_10_529 VPWR VGND sg13g2_fill_2
X_5677_ _2386_ net957 net774 VPWR VGND sg13g2_nand2_1
X_4628_ _1443_ _1440_ _1442_ VPWR VGND sg13g2_nand2_1
X_4559_ net834 net830 net880 net878 _1376_ VPWR VGND sg13g2_and4_1
X_6229_ net1051 VGND VPWR net182 mac2.sum_lvl2_ff\[40\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_18_618 VPWR VGND sg13g2_decap_8
XFILLER_46_938 VPWR VGND sg13g2_decap_8
XFILLER_17_139 VPWR VGND sg13g2_fill_1
XFILLER_25_161 VPWR VGND sg13g2_fill_1
XFILLER_13_345 VPWR VGND sg13g2_fill_1
XFILLER_40_131 VPWR VGND sg13g2_decap_4
XFILLER_1_750 VPWR VGND sg13g2_fill_2
XFILLER_37_916 VPWR VGND sg13g2_decap_8
X_3930_ _0775_ net1008 net922 net960 net920 VPWR VGND sg13g2_a22oi_1
XFILLER_45_993 VPWR VGND sg13g2_decap_8
XFILLER_16_183 VPWR VGND sg13g2_fill_1
X_3861_ _0705_ _0704_ _0687_ _0708_ VPWR VGND sg13g2_a21o_1
X_3792_ _0641_ net973 net916 VPWR VGND sg13g2_nand2_1
XFILLER_13_890 VPWR VGND sg13g2_fill_2
X_5600_ mac1.total_sum\[6\] mac2.total_sum\[6\] _2320_ VPWR VGND sg13g2_and2_1
XFILLER_9_850 VPWR VGND sg13g2_fill_1
X_5531_ VPWR VGND _2261_ _2260_ _2259_ mac2.sum_lvl3_ff\[25\] _2267_ net418 sg13g2_a221oi_1
XFILLER_8_371 VPWR VGND sg13g2_fill_1
X_5462_ net525 VPWR _2214_ VGND _2208_ _2212_ sg13g2_o21ai_1
X_5393_ _2160_ mac1.sum_lvl3_ff\[27\] mac1.sum_lvl3_ff\[7\] VPWR VGND sg13g2_nand2_1
X_4413_ _1239_ _1236_ _0128_ VPWR VGND sg13g2_xor2_1
XFILLER_28_1014 VPWR VGND sg13g2_decap_8
X_4344_ _1172_ _1122_ _1170_ VPWR VGND sg13g2_xnor2_1
X_6014_ net1078 VGND VPWR _0124_ mac1.products_ff\[75\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_4275_ _1094_ _1102_ _1104_ _1105_ VPWR VGND sg13g2_or3_1
X_3226_ _2816_ _2815_ _0104_ VPWR VGND sg13g2_xor2_1
XFILLER_28_916 VPWR VGND sg13g2_decap_8
XFILLER_39_220 VPWR VGND sg13g2_fill_1
X_3157_ _2744_ VPWR _2749_ VGND _2746_ _2747_ sg13g2_o21ai_1
X_3088_ _2679_ _2680_ _2674_ _2682_ VPWR VGND sg13g2_nand3_1
XFILLER_23_610 VPWR VGND sg13g2_fill_1
XFILLER_10_326 VPWR VGND sg13g2_fill_1
X_5729_ net926 net909 net775 _2437_ VPWR VGND sg13g2_mux2_1
Xheichips25_SDR_39 VPWR VGND uio_oe[6] sg13g2_tiehi
Xhold371 _0022_ VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold360 _2296_ VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold393 mac1.sum_lvl3_ff\[2\] VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold382 DP_2.matrix\[5\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xfanout840 net298 net840 VPWR VGND sg13g2_buf_8
Xfanout851 net302 net851 VPWR VGND sg13g2_buf_8
Xfanout873 net396 net873 VPWR VGND sg13g2_buf_8
Xfanout862 net497 net862 VPWR VGND sg13g2_buf_8
Xfanout884 net370 net884 VPWR VGND sg13g2_buf_8
XFILLER_45_201 VPWR VGND sg13g2_fill_1
Xfanout895 net301 net895 VPWR VGND sg13g2_buf_8
XFILLER_33_418 VPWR VGND sg13g2_fill_1
XFILLER_34_919 VPWR VGND sg13g2_decap_8
XFILLER_26_61 VPWR VGND sg13g2_fill_2
XFILLER_26_492 VPWR VGND sg13g2_fill_1
XFILLER_42_952 VPWR VGND sg13g2_decap_8
XFILLER_41_451 VPWR VGND sg13g2_fill_1
XFILLER_3_10 VPWR VGND sg13g2_fill_1
X_4060_ _0888_ _0883_ _0890_ _0901_ VPWR VGND sg13g2_a21o_1
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
X_3011_ _2604_ _2605_ _2607_ _2608_ VPWR VGND sg13g2_nor3_1
XFILLER_36_201 VPWR VGND sg13g2_fill_1
XFILLER_37_779 VPWR VGND sg13g2_fill_1
XFILLER_33_930 VPWR VGND sg13g2_decap_8
X_4962_ _1762_ _1761_ _1758_ VPWR VGND sg13g2_nand2b_1
X_4893_ _1674_ VPWR _1700_ VGND _1643_ _1672_ sg13g2_o21ai_1
X_3913_ _0758_ _0757_ _0754_ VPWR VGND sg13g2_nand2b_1
X_3844_ _0690_ _0657_ _0691_ VPWR VGND sg13g2_xor2_1
X_3775_ net924 net918 net973 net972 _0625_ VPWR VGND sg13g2_and4_1
X_6494_ net1031 VGND VPWR net14 DP_3.I_range.out_data\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5514_ mac2.sum_lvl3_ff\[22\] net451 _2254_ VPWR VGND sg13g2_and2_1
X_5445_ net321 _2198_ _0040_ VPWR VGND sg13g2_xor2_1
X_5376_ _2147_ mac1.sum_lvl3_ff\[23\] mac1.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
X_4327_ _1154_ _1153_ _1119_ _1156_ VPWR VGND sg13g2_a21o_1
X_4258_ _1088_ _1082_ _1086_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_1011 VPWR VGND sg13g2_decap_8
X_3209_ _2800_ net1006 net901 net942 net897 VPWR VGND sg13g2_a22oi_1
X_4189_ _1020_ _1002_ _0083_ VPWR VGND sg13g2_xor2_1
XFILLER_42_215 VPWR VGND sg13g2_fill_2
XFILLER_24_974 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_fill_1
XFILLER_7_606 VPWR VGND sg13g2_decap_8
Xhold190 mac1.products_ff\[7\] VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_46_510 VPWR VGND sg13g2_fill_2
XFILLER_18_201 VPWR VGND sg13g2_fill_2
XFILLER_46_532 VPWR VGND sg13g2_fill_1
XFILLER_46_554 VPWR VGND sg13g2_decap_8
XFILLER_46_587 VPWR VGND sg13g2_fill_2
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_30_955 VPWR VGND sg13g2_decap_8
XFILLER_41_292 VPWR VGND sg13g2_fill_1
X_3560_ _0419_ _0420_ _0385_ _0421_ VPWR VGND sg13g2_nand3_1
XFILLER_6_650 VPWR VGND sg13g2_fill_2
X_5230_ _2021_ _2010_ _2023_ VPWR VGND sg13g2_xor2_1
X_3491_ _0353_ _0347_ _0351_ VPWR VGND sg13g2_xnor2_1
X_5161_ _1956_ net844 net785 VPWR VGND sg13g2_nand2_1
X_4112_ _0949_ _0932_ _0952_ VPWR VGND sg13g2_xor2_1
X_5092_ _1865_ _1886_ _1888_ _1889_ VPWR VGND sg13g2_or3_1
X_4043_ _0885_ net966 net908 VPWR VGND sg13g2_nand2_2
XFILLER_25_716 VPWR VGND sg13g2_fill_1
X_5994_ net1064 VGND VPWR _0072_ mac1.products_ff\[3\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_4945_ _1746_ net847 net799 net849 net795 VPWR VGND sg13g2_a22oi_1
XFILLER_33_29 VPWR VGND sg13g2_fill_1
X_4876_ _1682_ _1668_ _1684_ VPWR VGND sg13g2_xor2_1
XFILLER_21_955 VPWR VGND sg13g2_decap_8
X_3827_ _0673_ _0672_ _0655_ _0675_ VPWR VGND sg13g2_a21o_1
X_3758_ _0612_ _0598_ _0611_ VPWR VGND sg13g2_xnor2_1
X_6477_ net1013 VGND VPWR net420 mac2.total_sum\[5\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3689_ _0545_ _0519_ _0546_ VPWR VGND sg13g2_xor2_1
X_5428_ _2188_ mac1.sum_lvl3_ff\[34\] net373 VPWR VGND sg13g2_nand2_1
XFILLER_0_848 VPWR VGND sg13g2_fill_2
X_5359_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] _2135_ VPWR VGND sg13g2_nor2_1
XFILLER_28_510 VPWR VGND sg13g2_fill_2
XFILLER_28_565 VPWR VGND sg13g2_decap_8
XFILLER_16_727 VPWR VGND sg13g2_fill_2
XFILLER_15_248 VPWR VGND sg13g2_decap_4
XFILLER_12_999 VPWR VGND sg13g2_decap_8
XFILLER_8_959 VPWR VGND sg13g2_decap_8
XFILLER_48_1017 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_686 VPWR VGND sg13g2_fill_1
XFILLER_24_8 VPWR VGND sg13g2_fill_1
XFILLER_34_568 VPWR VGND sg13g2_fill_2
X_2991_ VPWR _2591_ net1005 VGND sg13g2_inv_1
X_4730_ _1541_ _1533_ _1542_ VPWR VGND sg13g2_nor2b_1
X_4661_ _1472_ _1473_ _1456_ _1475_ VPWR VGND sg13g2_nand3_1
X_6400_ net1093 VGND VPWR net261 mac2.sum_lvl1_ff\[13\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3612_ _0439_ _0433_ _0441_ _0471_ VPWR VGND sg13g2_a21o_1
X_6331_ net1016 VGND VPWR net408 mac1.total_sum\[8\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_4592_ _1406_ _1407_ _1389_ _1408_ VPWR VGND sg13g2_nand3_1
XFILLER_7_992 VPWR VGND sg13g2_decap_8
X_3543_ _0364_ VPWR _0404_ VGND _0362_ _0365_ sg13g2_o21ai_1
X_3474_ _0335_ _0334_ _0325_ _0337_ VPWR VGND sg13g2_a21o_1
X_6262_ net1051 VGND VPWR net234 mac2.sum_lvl1_ff\[75\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5213_ _1994_ VPWR _2006_ VGND _1986_ _1995_ sg13g2_o21ai_1
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
X_6193_ net1096 VGND VPWR net103 mac1.sum_lvl2_ff\[14\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5144_ _1940_ _1896_ _1899_ VPWR VGND sg13g2_nand2_1
X_5075_ _1872_ _1826_ _1869_ VPWR VGND sg13g2_xnor2_1
X_4026_ _0867_ _0868_ _0869_ VPWR VGND sg13g2_nor2b_1
X_5977_ net801 _0259_ VPWR VGND sg13g2_buf_1
X_4928_ _1726_ _1727_ _1729_ _1730_ VPWR VGND sg13g2_nor3_1
X_4859_ _1655_ VPWR _1667_ VGND _1635_ _1656_ sg13g2_o21ai_1
XFILLER_0_634 VPWR VGND sg13g2_fill_2
XFILLER_29_874 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_fill_1
XFILLER_7_200 VPWR VGND sg13g2_fill_1
XFILLER_4_940 VPWR VGND sg13g2_decap_8
X_3190_ _2781_ net957 net1003 VPWR VGND sg13g2_nand2_1
X_5900_ _2578_ net825 net759 VPWR VGND sg13g2_nand2_1
XFILLER_46_170 VPWR VGND sg13g2_fill_2
XFILLER_35_866 VPWR VGND sg13g2_decap_8
X_5831_ VGND VPWR net754 _2533_ _0174_ _2531_ sg13g2_a21oi_1
X_5762_ net867 net882 net780 _2469_ VPWR VGND sg13g2_mux2_1
X_4713_ _1479_ VPWR _1526_ VGND _1419_ _1480_ sg13g2_o21ai_1
X_5693_ net981 DP_1.matrix\[42\] net775 _2402_ VPWR VGND sg13g2_mux2_1
X_4644_ _1458_ net826 net879 VPWR VGND sg13g2_nand2_1
X_4575_ _1391_ net883 net823 VPWR VGND sg13g2_nand2_1
X_3526_ _0387_ DP_1.matrix\[0\] net1005 VPWR VGND sg13g2_nand2_1
X_6314_ net1036 VGND VPWR net67 mac2.sum_lvl3_ff\[27\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6245_ net1039 VGND VPWR net249 mac1.sum_lvl1_ff\[74\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3457_ _0320_ net991 net927 VPWR VGND sg13g2_nand2_1
X_3388_ _2969_ net358 net929 VPWR VGND sg13g2_nand2_1
X_6176_ net1083 VGND VPWR net210 mac1.sum_lvl1_ff\[49\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_5127_ net794 net791 net839 net997 _1923_ VPWR VGND sg13g2_and4_1
X_5058_ _1844_ VPWR _1855_ VGND _1823_ _1845_ sg13g2_o21ai_1
X_4009_ _0852_ net966 net910 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_64_clk clknet_4_2_0_clk clknet_leaf_64_clk VPWR VGND sg13g2_buf_8
XFILLER_26_866 VPWR VGND sg13g2_decap_8
XFILLER_38_1005 VPWR VGND sg13g2_decap_8
XFILLER_4_236 VPWR VGND sg13g2_fill_1
XFILLER_1_976 VPWR VGND sg13g2_decap_8
XFILLER_49_947 VPWR VGND sg13g2_decap_8
Xhold50 mac2.sum_lvl1_ff\[4\] VPWR VGND net90 sg13g2_dlygate4sd3_1
Xhold61 mac1.sum_lvl1_ff\[4\] VPWR VGND net101 sg13g2_dlygate4sd3_1
Xhold83 mac1.sum_lvl2_ff\[48\] VPWR VGND net123 sg13g2_dlygate4sd3_1
Xhold72 mac2.products_ff\[79\] VPWR VGND net112 sg13g2_dlygate4sd3_1
Xhold94 mac1.products_ff\[71\] VPWR VGND net134 sg13g2_dlygate4sd3_1
XFILLER_44_641 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_55_clk clknet_4_8_0_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
XFILLER_6_10 VPWR VGND sg13g2_fill_1
X_4360_ _1186_ _1187_ _1188_ VPWR VGND sg13g2_nor2_1
X_3311_ _2897_ _2886_ _2899_ VPWR VGND sg13g2_xor2_1
X_4291_ _1092_ VPWR _1120_ VGND _1090_ _1093_ sg13g2_o21ai_1
X_6030_ net1076 VGND VPWR _0167_ DP_3.matrix\[44\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_6_1003 VPWR VGND sg13g2_decap_8
X_3242_ _2832_ net947 net890 VPWR VGND sg13g2_nand2_1
X_3173_ VGND VPWR _2761_ _2762_ _2765_ _2743_ sg13g2_a21oi_1
Xfanout1092 net1095 net1092 VPWR VGND sg13g2_buf_8
Xfanout1081 net1082 net1081 VPWR VGND sg13g2_buf_8
Xfanout1070 net1071 net1070 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_46_clk clknet_4_14_0_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
X_5814_ _2517_ VPWR _2520_ VGND _2518_ _2519_ sg13g2_o21ai_1
X_5745_ DP_3.Q_range.out_data\[2\] _2589_ DP_3.Q_range.out_data\[4\] DP_3.Q_range.out_data\[6\]
+ _2452_ VPWR VGND sg13g2_nor4_1
X_5676_ net991 net776 _2385_ VPWR VGND sg13g2_nor2_1
X_4627_ _1439_ _1438_ _1421_ _1442_ VPWR VGND sg13g2_a21o_1
X_4558_ _1375_ net883 net827 VPWR VGND sg13g2_nand2_1
X_4489_ _1313_ _1312_ _1285_ VPWR VGND sg13g2_nand2b_1
X_3509_ _0360_ _0368_ _0370_ _0371_ VPWR VGND sg13g2_or3_1
X_6228_ net1052 VGND VPWR net235 mac2.sum_lvl2_ff\[39\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6159_ net1060 VGND VPWR _0264_ DP_4.matrix\[76\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_46_917 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_37_clk clknet_4_14_0_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_26_696 VPWR VGND sg13g2_decap_8
XFILLER_40_165 VPWR VGND sg13g2_decap_4
XFILLER_1_762 VPWR VGND sg13g2_fill_1
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_36_405 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_28_clk clknet_4_6_0_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_36_449 VPWR VGND sg13g2_fill_2
XFILLER_45_972 VPWR VGND sg13g2_decap_8
XFILLER_32_611 VPWR VGND sg13g2_fill_1
X_3860_ VGND VPWR _0704_ _0705_ _0707_ _0687_ sg13g2_a21oi_1
X_3791_ _0626_ VPWR _0640_ VGND _0624_ _0627_ sg13g2_o21ai_1
XFILLER_9_862 VPWR VGND sg13g2_fill_1
XFILLER_9_840 VPWR VGND sg13g2_fill_1
X_5530_ _2266_ mac2.sum_lvl3_ff\[26\] net457 VPWR VGND sg13g2_xnor2_1
XFILLER_31_187 VPWR VGND sg13g2_fill_1
XFILLER_9_873 VPWR VGND sg13g2_fill_1
X_5461_ _2208_ net525 _2212_ _2213_ VPWR VGND sg13g2_nor3_2
X_4412_ _1239_ _1237_ _1238_ VPWR VGND sg13g2_nand2b_1
X_5392_ _2158_ net485 _0028_ VPWR VGND sg13g2_nor2b_1
X_4343_ VGND VPWR _1171_ _1169_ _1123_ sg13g2_or2_1
X_4274_ VGND VPWR _1100_ _1101_ _1104_ _1095_ sg13g2_a21oi_1
X_6013_ net1068 VGND VPWR _0123_ mac1.products_ff\[74\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3225_ _2816_ _2773_ _2776_ VPWR VGND sg13g2_nand2_1
X_3156_ _2744_ _2746_ _2747_ _2748_ VPWR VGND sg13g2_nor3_1
X_3087_ _2681_ _2674_ _2679_ _2680_ VPWR VGND sg13g2_and3_1
Xclkbuf_leaf_19_clk clknet_4_4_0_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_36_983 VPWR VGND sg13g2_decap_8
X_5728_ _2413_ _2435_ _2436_ VPWR VGND sg13g2_nor2b_1
X_3989_ _0791_ _0788_ _0831_ _0833_ VPWR VGND sg13g2_a21o_1
X_5659_ _2359_ _2362_ _2368_ VPWR VGND sg13g2_nor2_1
Xhold350 DP_2.matrix\[44\] VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold361 _0052_ VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold372 DP_1.matrix\[37\] VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold394 _2145_ VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold383 mac2.sum_lvl3_ff\[31\] VPWR VGND net423 sg13g2_dlygate4sd3_1
Xfanout841 net843 net841 VPWR VGND sg13g2_buf_8
Xfanout852 DP_3.matrix\[73\] net852 VPWR VGND sg13g2_buf_8
Xfanout830 DP_4.matrix\[1\] net830 VPWR VGND sg13g2_buf_1
Xfanout874 net386 net874 VPWR VGND sg13g2_buf_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
Xfanout885 DP_3.matrix\[1\] net885 VPWR VGND sg13g2_buf_1
Xfanout863 net864 net863 VPWR VGND sg13g2_buf_8
Xfanout896 net897 net896 VPWR VGND sg13g2_buf_8
XFILLER_46_736 VPWR VGND sg13g2_fill_1
XFILLER_42_931 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_fill_1
X_3010_ _2607_ net952 net903 net954 net899 VPWR VGND sg13g2_a22oi_1
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_983 VPWR VGND sg13g2_decap_8
X_4961_ _1760_ _1739_ _1761_ VPWR VGND sg13g2_xor2_1
X_4892_ _1699_ _1694_ _1697_ VPWR VGND sg13g2_xnor2_1
X_3912_ _0756_ _0717_ _0757_ VPWR VGND sg13g2_xor2_1
X_3843_ _0690_ net972 net914 VPWR VGND sg13g2_nand2_1
XFILLER_20_625 VPWR VGND sg13g2_fill_2
XFILLER_32_474 VPWR VGND sg13g2_fill_2
XFILLER_33_986 VPWR VGND sg13g2_decap_8
X_3774_ _0624_ net975 net916 VPWR VGND sg13g2_nand2_1
X_6493_ net1031 VGND VPWR net13 DP_3.I_range.out_data\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_5513_ _2250_ VPWR _2253_ VGND _2249_ _2251_ sg13g2_o21ai_1
Xclkbuf_leaf_8_clk clknet_4_3_0_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5444_ net320 mac2.sum_lvl2_ff\[21\] _2200_ VPWR VGND sg13g2_xor2_1
X_5375_ VGND VPWR _2144_ _2146_ _2145_ _2143_ sg13g2_a21oi_2
X_4326_ _1153_ _1154_ _1119_ _1155_ VPWR VGND sg13g2_nand3_1
X_4257_ _1082_ _1086_ _1087_ VPWR VGND sg13g2_and2_1
X_3208_ net901 net897 net941 net1006 _2799_ VPWR VGND sg13g2_and4_1
X_4188_ _1002_ _1020_ _1021_ VPWR VGND sg13g2_and2_1
XFILLER_28_725 VPWR VGND sg13g2_fill_1
X_3139_ _2730_ _2729_ _0102_ VPWR VGND sg13g2_xor2_1
XFILLER_43_706 VPWR VGND sg13g2_fill_2
XFILLER_24_953 VPWR VGND sg13g2_decap_8
XFILLER_6_139 VPWR VGND sg13g2_fill_2
XFILLER_3_824 VPWR VGND sg13g2_fill_1
Xhold180 mac1.sum_lvl1_ff\[48\] VPWR VGND net220 sg13g2_dlygate4sd3_1
Xhold191 mac1.products_ff\[70\] VPWR VGND net231 sg13g2_dlygate4sd3_1
XFILLER_46_500 VPWR VGND sg13g2_fill_1
XFILLER_34_706 VPWR VGND sg13g2_fill_1
XFILLER_14_452 VPWR VGND sg13g2_fill_1
XFILLER_14_463 VPWR VGND sg13g2_fill_1
XFILLER_18_1025 VPWR VGND sg13g2_decap_4
XFILLER_30_934 VPWR VGND sg13g2_decap_8
X_3490_ _0347_ _0351_ _0352_ VPWR VGND sg13g2_and2_1
X_5160_ VGND VPWR net794 net838 _1955_ _1922_ sg13g2_a21oi_1
X_4111_ _0932_ _0949_ _0951_ VPWR VGND sg13g2_nor2_1
X_5091_ VGND VPWR _1884_ _1885_ _1888_ _1866_ sg13g2_a21oi_1
X_4042_ _0884_ net971 net1004 VPWR VGND sg13g2_nand2_1
X_5993_ net1045 VGND VPWR _0071_ mac1.products_ff\[2\] clknet_leaf_55_clk sg13g2_dfrbpq_1
XFILLER_18_791 VPWR VGND sg13g2_fill_1
X_4944_ net795 net849 net799 _1745_ VPWR VGND net847 sg13g2_nand4_1
X_4875_ _1683_ _1668_ _1682_ VPWR VGND sg13g2_nand2_1
XFILLER_20_411 VPWR VGND sg13g2_fill_2
XFILLER_21_934 VPWR VGND sg13g2_decap_8
X_3826_ _0672_ _0673_ _0655_ _0674_ VPWR VGND sg13g2_nand3_1
X_3757_ _0611_ _0608_ _0610_ VPWR VGND sg13g2_xnor2_1
X_6476_ net1013 VGND VPWR net456 mac2.total_sum\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3688_ _0545_ net982 DP_2.matrix\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_0_805 VPWR VGND sg13g2_fill_2
X_5427_ _0020_ _2184_ net342 VPWR VGND sg13g2_xnor2_1
XFILLER_0_838 VPWR VGND sg13g2_fill_1
X_5358_ _2134_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
X_4309_ _1098_ VPWR _1138_ VGND _1096_ _1099_ sg13g2_o21ai_1
X_5289_ _2079_ net838 net994 VPWR VGND sg13g2_nand2_1
XFILLER_15_205 VPWR VGND sg13g2_fill_1
XFILLER_43_547 VPWR VGND sg13g2_fill_1
XFILLER_8_938 VPWR VGND sg13g2_decap_8
XFILLER_7_404 VPWR VGND sg13g2_fill_1
XFILLER_12_978 VPWR VGND sg13g2_decap_8
XFILLER_23_293 VPWR VGND sg13g2_fill_2
XFILLER_7_426 VPWR VGND sg13g2_fill_2
XFILLER_11_499 VPWR VGND sg13g2_fill_1
XFILLER_3_0 VPWR VGND sg13g2_fill_1
XFILLER_19_544 VPWR VGND sg13g2_fill_1
XFILLER_19_555 VPWR VGND sg13g2_fill_2
XFILLER_47_897 VPWR VGND sg13g2_decap_8
X_2990_ VPWR _2590_ net1010 VGND sg13g2_inv_1
X_4660_ _1474_ _1456_ _1472_ _1473_ VPWR VGND sg13g2_and3_1
X_3611_ _0470_ _0469_ _0115_ VPWR VGND sg13g2_xor2_1
XFILLER_31_1011 VPWR VGND sg13g2_decap_8
XFILLER_7_971 VPWR VGND sg13g2_decap_8
X_6330_ net1013 VGND VPWR net521 mac1.total_sum\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4591_ _1395_ VPWR _1407_ VGND _1403_ _1405_ sg13g2_o21ai_1
X_3542_ _0403_ _0397_ _0402_ VPWR VGND sg13g2_xnor2_1
X_3473_ _0334_ _0335_ _0325_ _0336_ VPWR VGND sg13g2_nand3_1
X_6261_ net1052 VGND VPWR net252 mac2.sum_lvl1_ff\[74\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
X_6192_ net1085 VGND VPWR net110 mac1.sum_lvl2_ff\[13\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5212_ _0151_ _2004_ _2005_ VPWR VGND sg13g2_xnor2_1
X_5143_ _1936_ _1938_ _1939_ VPWR VGND sg13g2_nor2_1
X_5074_ _1826_ _1869_ _1871_ VPWR VGND sg13g2_and2_1
XFILLER_49_190 VPWR VGND sg13g2_fill_1
X_4025_ _0830_ _0866_ _0828_ _0868_ VPWR VGND sg13g2_nand3_1
XFILLER_25_503 VPWR VGND sg13g2_fill_2
XFILLER_38_886 VPWR VGND sg13g2_decap_8
X_5976_ net803 _0258_ VPWR VGND sg13g2_buf_1
XFILLER_12_208 VPWR VGND sg13g2_fill_1
X_4927_ _1729_ net849 net799 net850 DP_4.matrix\[73\] VPWR VGND sg13g2_a22oi_1
X_4858_ _1665_ _1661_ _0141_ VPWR VGND sg13g2_xor2_1
X_3809_ _0657_ net974 net912 VPWR VGND sg13g2_nand2_1
XFILLER_20_252 VPWR VGND sg13g2_fill_1
XFILLER_21_797 VPWR VGND sg13g2_fill_2
XFILLER_5_908 VPWR VGND sg13g2_fill_2
X_4789_ _1600_ _1571_ _1598_ VPWR VGND sg13g2_xnor2_1
X_6459_ net1062 VGND VPWR net362 mac2.sum_lvl3_ff\[3\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_47_127 VPWR VGND sg13g2_fill_1
XFILLER_18_52 VPWR VGND sg13g2_fill_2
XFILLER_24_580 VPWR VGND sg13g2_fill_1
XFILLER_11_241 VPWR VGND sg13g2_fill_2
XFILLER_8_768 VPWR VGND sg13g2_fill_1
XFILLER_4_996 VPWR VGND sg13g2_decap_8
XFILLER_38_138 VPWR VGND sg13g2_fill_2
X_5830_ _2533_ _2394_ _2532_ VPWR VGND sg13g2_nand2_1
XFILLER_34_366 VPWR VGND sg13g2_fill_1
X_5761_ _2462_ _2467_ _2468_ VPWR VGND sg13g2_nor2b_1
X_4712_ _1522_ _1523_ _1454_ _1525_ VPWR VGND sg13g2_nand3_1
X_5692_ _2378_ _2400_ _2401_ VPWR VGND sg13g2_nor2b_1
X_4643_ _1457_ net883 net822 VPWR VGND sg13g2_nand2_1
X_4574_ _1390_ net886 net822 VPWR VGND sg13g2_nand2_1
X_3525_ _0358_ VPWR _0386_ VGND _0355_ _0359_ sg13g2_o21ai_1
X_6313_ net1036 VGND VPWR net117 mac2.sum_lvl3_ff\[26\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6244_ net1040 VGND VPWR net51 mac1.sum_lvl1_ff\[73\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3456_ _0302_ VPWR _0319_ VGND _0293_ _0303_ sg13g2_o21ai_1
X_3387_ _2967_ _2961_ _0071_ VPWR VGND sg13g2_xor2_1
X_6175_ net1083 VGND VPWR net232 mac1.sum_lvl1_ff\[48\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5126_ _1922_ net791 net998 VPWR VGND sg13g2_nand2_1
X_5057_ _1853_ _1852_ _0157_ VPWR VGND sg13g2_xor2_1
X_4008_ VGND VPWR net919 net960 _0851_ _0818_ sg13g2_a21oi_1
XFILLER_26_845 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
X_5959_ net861 _0233_ VPWR VGND sg13g2_buf_1
XFILLER_4_204 VPWR VGND sg13g2_fill_2
XFILLER_5_749 VPWR VGND sg13g2_fill_1
XFILLER_49_926 VPWR VGND sg13g2_decap_8
XFILLER_1_955 VPWR VGND sg13g2_decap_8
Xhold40 mac1.products_ff\[15\] VPWR VGND net80 sg13g2_dlygate4sd3_1
Xhold62 mac1.products_ff\[151\] VPWR VGND net102 sg13g2_dlygate4sd3_1
Xhold73 mac2.sum_lvl2_ff\[47\] VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold51 mac2.sum_lvl1_ff\[86\] VPWR VGND net91 sg13g2_dlygate4sd3_1
Xhold84 mac2.sum_lvl1_ff\[15\] VPWR VGND net124 sg13g2_dlygate4sd3_1
Xhold95 mac1.sum_lvl1_ff\[10\] VPWR VGND net135 sg13g2_dlygate4sd3_1
XFILLER_16_311 VPWR VGND sg13g2_fill_2
XFILLER_40_892 VPWR VGND sg13g2_decap_8
XFILLER_8_576 VPWR VGND sg13g2_fill_1
X_3310_ VGND VPWR _2898_ _2897_ _2886_ sg13g2_or2_1
X_4290_ _1108_ VPWR _1119_ VGND _1088_ _1109_ sg13g2_o21ai_1
X_3241_ VGND VPWR net901 net942 _2831_ _2798_ sg13g2_a21oi_1
X_3172_ _2761_ _2762_ _2743_ _2764_ VPWR VGND sg13g2_nand3_1
Xfanout1082 net1087 net1082 VPWR VGND sg13g2_buf_8
Xfanout1071 net1077 net1071 VPWR VGND sg13g2_buf_8
Xfanout1060 net1062 net1060 VPWR VGND sg13g2_buf_8
Xfanout1093 net1094 net1093 VPWR VGND sg13g2_buf_8
XFILLER_19_193 VPWR VGND sg13g2_decap_4
X_5813_ net768 VPWR _2519_ VGND net821 net778 sg13g2_o21ai_1
XFILLER_34_174 VPWR VGND sg13g2_decap_4
X_5744_ VGND VPWR _2592_ net777 _2451_ _2450_ sg13g2_a21oi_1
X_5675_ _2384_ net770 _2383_ net763 net959 VPWR VGND sg13g2_a22oi_1
XFILLER_31_892 VPWR VGND sg13g2_decap_8
X_4626_ VGND VPWR _1438_ _1439_ _1441_ _1421_ sg13g2_a21oi_1
X_4557_ _1360_ VPWR _1374_ VGND _1358_ _1361_ sg13g2_o21ai_1
X_4488_ _1310_ _1271_ _1312_ VPWR VGND sg13g2_xor2_1
X_3508_ VGND VPWR _0366_ _0367_ _0370_ _0361_ sg13g2_a21oi_1
X_3439_ VGND VPWR _0299_ _0300_ _0303_ _0294_ sg13g2_a21oi_1
X_6227_ net1052 VGND VPWR net196 mac2.sum_lvl2_ff\[38\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6158_ net1054 VGND VPWR _0263_ DP_4.matrix\[75\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_5109_ _1905_ net848 net781 VPWR VGND sg13g2_nand2_1
X_6089_ net1042 VGND VPWR _0212_ DP_2.matrix\[72\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_25_130 VPWR VGND sg13g2_fill_2
XFILLER_25_152 VPWR VGND sg13g2_fill_2
XFILLER_15_97 VPWR VGND sg13g2_fill_1
XFILLER_40_199 VPWR VGND sg13g2_decap_4
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_49_778 VPWR VGND sg13g2_decap_8
XFILLER_45_951 VPWR VGND sg13g2_decap_8
XFILLER_17_653 VPWR VGND sg13g2_fill_1
X_3790_ VGND VPWR _0639_ _0638_ _0636_ sg13g2_or2_1
XFILLER_32_678 VPWR VGND sg13g2_fill_2
XFILLER_13_892 VPWR VGND sg13g2_fill_1
X_5460_ VPWR VGND _2206_ _2205_ _2204_ mac2.sum_lvl2_ff\[24\] _2212_ mac2.sum_lvl2_ff\[5\]
+ sg13g2_a221oi_1
X_4411_ VGND VPWR _1160_ _1200_ _1238_ _1201_ sg13g2_a21oi_1
X_5391_ net484 VPWR _2159_ VGND _2153_ _2157_ sg13g2_o21ai_1
X_4342_ _1170_ net866 net804 VPWR VGND sg13g2_nand2_1
X_4273_ _1100_ _1101_ _1095_ _1103_ VPWR VGND sg13g2_nand3_1
X_6012_ net1068 VGND VPWR _0116_ mac1.products_ff\[73\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3224_ _2812_ _2814_ _2815_ VPWR VGND sg13g2_nor2_1
.ends

